//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "MUX2.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [7:0] w3;    //: /sn:0 {0}(#:220,76)(220,92){1}
//: {2}(#:218,94)(110,94)(110,70){3}
//: {4}(220,96)(220,109){5}
reg [7:0] w1;    //: /sn:0 {0}(#:332,77)(332,92){1}
//: {2}(#:334,94)(449,94)(449,71){3}
//: {4}(332,96)(332,109){5}
reg w2;    //: /sn:0 {0}(427,135)(381,135){1}
reg w10;    //: /sn:0 {0}(82,181)(179,181){1}
reg w9;    //: /sn:0 {0}(82,132)(179,132){1}
wire [8:0] w6;    //: /sn:0 {0}(#:157,255)(175,255){1}
//: {2}(179,255)(222,255)(#:222,220){3}
//: {4}(#:177,257)(177,293)(158,293){5}
wire [7:0] w7;    //: /sn:0 {0}(#:351,220)(351,244)(352,244){1}
//: {2}(356,244)(390,244){3}
//: {4}(#:354,246)(354,276)(370,276){5}
wire [7:0] w8;    //: /sn:0 {0}(#:449,182)(449,191)(435,191){1}
//: {2}(431,191)(#:381,191){3}
//: {4}(#:433,193)(433,208)(452,208){5}
wire [15:0] w5;    //: /sn:0 {0}(#:284,269)(286,269)(286,256){1}
//: {2}(#:288,254)(318,254)(318,306)(295,306){3}
//: {4}(286,252)(#:286,220){5}
//: enddecls

  //: LED g4 (w8) @(449,175) /sn:0 /w:[ 0 ] /type:1
  //: LED g8 (w6) @(151,293) /sn:0 /R:1 /w:[ 5 ] /type:3
  //: SWITCH g3 (w2) @(445,135) /sn:0 /R:2 /w:[ 0 ] /st:0 /dn:1
  //: LED g13 (w7) @(397,244) /sn:0 /R:3 /w:[ 3 ] /type:1
  //: SWITCH g2 (w10) @(65,181) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g1 (w9) @(65,132) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g11 (w5) @(288,306) /sn:0 /R:1 /w:[ 3 ] /type:3
  //: LED g16 (w8) @(459,208) /sn:0 /R:3 /w:[ 5 ] /type:3
  //: LED g10 (w5) @(277,269) /sn:0 /R:1 /w:[ 0 ] /type:1
  //: joint g19 (w3) @(220, 94) /w:[ -1 1 2 4 ]
  //: DIP g6 (w1) @(332,67) /sn:0 /w:[ 0 ] /st:3 /dn:1
  //: LED g7 (w6) @(150,255) /sn:0 /R:1 /w:[ 0 ] /type:1
  //: joint g9 (w6) @(177, 255) /w:[ 2 -1 1 4 ]
  //: joint g15 (w7) @(354, 244) /w:[ 2 -1 1 4 ]
  //: LED g20 (w1) @(449,64) /sn:0 /w:[ 3 ] /type:3
  //: joint g17 (w8) @(433, 191) /w:[ 1 -1 2 4 ]
  //: DIP g5 (w3) @(220,66) /sn:0 /w:[ 0 ] /st:9 /dn:1
  //: LED g14 (w7) @(377,276) /sn:0 /R:3 /w:[ 5 ] /type:3
  //: joint g21 (w1) @(332, 94) /w:[ 2 1 -1 4 ]
  Calcolatrice_4_operazioni g0 (.A(w3), .B(w1), .Neg(w10), .Clk(w9), .Carica(w2), .AdivB(w7), .AddSub(w6), .AxB(w5), .RestoDiv(w8));   //: @(180, 110) /sz:(200, 109) /sn:0 /p:[ Ti0>5 Ti1>5 Li0>1 Li1>1 Ri0>1 Bo0<0 Bo1<3 Bo2<5 Ro0<3 ]
  //: joint g12 (w5) @(286, 254) /w:[ 2 4 -1 1 ]
  //: LED g18 (w3) @(110,63) /sn:0 /w:[ 3 ] /type:3

endmodule
//: /netlistEnd

//: /netlistBegin NAND2
module NAND2(in1, out, in2);
//: interface  /sz:(40, 40) /bd:[ Li0>in1(10/40) Li1>in2(30/40) Ro0<out(18/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w6;    //: /sn:0 {0}(154,1)(154,4)(154,4)(154,13){1}
//: {2}(156,15)(182,15)(182,25){3}
//: {4}(152,15)(127,15)(127,42){5}
output out;    //: /sn:0 {0}(155,109)(155,90){1}
//: {2}(157,88)(169,88)(169,88)(218,88){3}
//: {4}(155,86)(155,76){5}
//: {6}(157,74)(182,74)(182,42){7}
//: {8}(153,74)(127,74)(127,59){9}
supply0 w3;    //: /sn:0 {0}(155,184)(155,208){1}
input in1;    //: /sn:0 {0}(46,33)(58,33)(58,33)(70,33){1}
//: {2}(74,33)(155,33)(155,33)(168,33){3}
//: {4}(72,35)(72,117)(141,117){5}
input in2;    //: /sn:0 {0}(47,125)(86,125)(86,125)(101,125){1}
//: {2}(103,123)(103,50)(113,50){3}
//: {4}(103,127)(103,175)(141,175){5}
wire w4;    //: /sn:0 {0}(155,126)(155,167){1}
//: enddecls

  //: IN g8 (in1) @(44,33) /sn:0 /w:[ 0 ]
  //: joint g4 (out) @(155, 74) /w:[ 6 -1 8 5 ]
  //: joint g13 (in2) @(103, 125) /w:[ -1 2 1 4 ]
  _GGNMOS #(2, 1) g3 (.Z(w4), .S(w3), .G(in2));   //: @(149,175) /sn:0 /w:[ 1 0 5 ]
  _GGPMOS #(2, 1) g2 (.Z(out), .S(w6), .G(in1));   //: @(176,33) /sn:0 /w:[ 7 3 3 ]
  _GGNMOS #(2, 1) g1 (.Z(out), .S(w4), .G(in1));   //: @(149,117) /sn:0 /w:[ 0 0 5 ]
  //: joint g11 (out) @(155, 88) /w:[ 2 4 -1 1 ]
  //: OUT g10 (out) @(215,88) /sn:0 /w:[ 3 ]
  //: VDD g6 (w6) @(165,1) /sn:0 /w:[ 0 ]
  //: IN g9 (in2) @(45,125) /sn:0 /w:[ 0 ]
  //: joint g7 (w6) @(154, 15) /w:[ 2 1 4 -1 ]
  //: GROUND g5 (w3) @(155,214) /sn:0 /w:[ 1 ]
  _GGPMOS #(2, 1) g0 (.Z(out), .S(w6), .G(in2));   //: @(121,50) /sn:0 /w:[ 9 5 3 ]
  //: joint g12 (in1) @(72, 33) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFSR
module FFSR(S, Y, clk, R);
//: interface  /sz:(40, 40) /bd:[ Li0>R(28/40) Li1>S(7/40) Bi0>clk(17/40) Ro0<Y(18/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input R;    //: /sn:0 {0}(300,174)(225,174)(225,201)(210,201){1}
input clk;    //: /sn:0 {0}(300,194)(267,194){1}
//: {2}(265,192)(265,127)(301,127){3}
//: {4}(265,196)(265,289){5}
input S;    //: /sn:0 {0}(214,102)(286,102)(286,107)(301,107){1}
output Y;    //: /sn:0 {0}(479,175)(508,175)(508,173)(523,173){1}
wire w0;    //: /sn:0 {0}(342,183)(381,183)(381,175)(396,175){1}
wire w3;    //: /sn:0 {0}(494,154)(479,154){1}
wire w1;    //: /sn:0 {0}(343,116)(381,116)(381,151)(396,151){1}
//: enddecls

  //: IN g4 (S) @(212,102) /sn:0 /w:[ 0 ]
  AND2 g3 (.in2(clk), .in1(S), .out(w1));   //: @(302, 97) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]
  AND2 g2 (.in2(clk), .in1(R), .out(w0));   //: @(301, 164) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  //: OUT g1 (Y) @(520,173) /sn:0 /w:[ 1 ]
  //: IN g6 (clk) @(265,291) /sn:0 /R:1 /w:[ 5 ]
  //: joint g7 (clk) @(265, 194) /w:[ 1 2 -1 4 ]
  //: IN g5 (R) @(208,201) /sn:0 /w:[ 1 ]
  LATCHSR g0 (.s(w1), .r(w0), .Y1(w3), .Y(Y));   //: @(397, 144) /sz:(81, 47) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mul16b
module Mul16b(B, A, S);
//: interface  /sz:(63, 64) /bd:[ Li0>B[7:0](44/64) Li1>A[7:0](16/64) Bo0<S[15:0](32/63) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] A;    //: /sn:0 {0}(#:613,67)(569,67){1}
//: {2}(568,67)(516,67){3}
//: {4}(515,67)(461,67){5}
//: {6}(460,67)(408,67){7}
//: {8}(407,67)(352,67){9}
//: {10}(351,67)(297,67){11}
//: {12}(296,67)(247,67){13}
//: {14}(246,67)(187,67){15}
//: {16}(186,67)(50,67){17}
//: {18}(49,67)(-3,67){19}
//: {20}(-4,67)(-59,67){21}
//: {22}(-60,67)(-112,67){23}
//: {24}(-113,67)(-164,67){25}
//: {26}(-165,67)(-217,67){27}
//: {28}(-218,67)(-270,67){29}
//: {30}(-271,67)(-299,67)(-299,67)(-326,67){31}
//: {32}(-327,67)(-413,67){33}
//: {34}(-414,67)(-464,67){35}
//: {36}(-465,67)(-519,67){37}
//: {38}(-520,67)(-574,67){39}
//: {40}(-575,67)(-626,67){41}
//: {42}(-627,67)(-684,67){43}
//: {44}(-685,67)(-739,67){45}
//: {46}(-740,67)(-793,67){47}
//: {48}(-794,67)(-877,67){49}
//: {50}(-878,67)(-928,67){51}
//: {52}(-929,67)(-986,67){53}
//: {54}(-987,67)(-1042,67){55}
//: {56}(-1043,67)(-1094,67){57}
//: {58}(-1095,67)(-1150,67){59}
//: {60}(-1151,67)(-1204,67){61}
//: {62}(-1205,67)(-1260,67){63}
//: {64}(-1261,67)(-1343,67){65}
//: {66}(-1344,67)(-1401,67){67}
//: {68}(-1402,67)(-1453,67){69}
//: {70}(-1454,67)(-1505,67){71}
//: {72}(-1506,67)(-1561,67){73}
//: {74}(-1562,67)(-1615,67){75}
//: {76}(-1616,67)(-1667,67){77}
//: {78}(-1668,67)(-1721,67){79}
//: {80}(-1722,67)(-1813,67){81}
//: {82}(-1814,67)(-1866,67){83}
//: {84}(-1867,67)(-1918,67){85}
//: {86}(-1919,67)(-1974,67){87}
//: {88}(-1975,67)(-2026,67){89}
//: {90}(-2027,67)(-2080,67){91}
//: {92}(-2081,67)(-2136,67){93}
//: {94}(-2137,67)(-2188,67){95}
//: {96}(-2189,67)(-2284,67){97}
//: {98}(-2285,67)(-2335,67){99}
//: {100}(-2336,67)(-2388,67){101}
//: {102}(-2389,67)(-2438,67){103}
//: {104}(-2439,67)(-2492,67){105}
//: {106}(-2493,67)(-2547,67){107}
//: {108}(-2548,67)(-2594,67){109}
//: {110}(-2595,67)(-2649,67){111}
//: {112}(-2650,67)(-2751,67){113}
//: {114}(-2752,67)(-2805,67){115}
//: {116}(-2806,67)(-2859,67){117}
//: {118}(-2860,67)(-2913,67){119}
//: {120}(-2914,67)(-2969,67){121}
//: {122}(-2970,67)(-3019,67){123}
//: {124}(-3020,67)(-3073,67){125}
//: {126}(-3074,67)(-3128,67){127}
//: {128}(-3129,67)(-3141,67){129}
output [15:0] S;    //: /sn:0 {0}(135,1867)(78,1867)(#:78,1803){1}
input [7:0] B;    //: /sn:0 {0}(#:615,98)(605,98)(605,98)(589,98){1}
//: {2}(588,98)(70,98){3}
//: {4}(69,98)(-392,98){5}
//: {6}(-393,98)(-857,98){7}
//: {8}(-858,98)(-1324,98){9}
//: {10}(-1325,98)(-1793,98){11}
//: {12}(-1794,98)(-2265,98){13}
//: {14}(-2266,98)(-2728,98){15}
//: {16}(-2729,98)(-2770,98){17}
wire w32;    //: /sn:0 {0}(-216,355)(-216,79)(-217,79)(-217,71){1}
wire w96;    //: /sn:0 {0}(-1961,399)(-1961,1090)(4,1090)(4,1158){1}
wire w73;    //: /sn:0 {0}(-1451,356)(-1451,79)(-1453,79)(-1453,71){1}
wire w45;    //: /sn:0 {0}(-560,396)(-560,642)(223,642)(223,678){1}
wire w160;    //: /sn:0 {0}(161,556)(161,662)(183,662)(183,677){1}
wire w214;    //: /sn:0 {0}(23,1216)(23,1305)(29,1305)(29,1320){1}
wire w203;    //: /sn:0 {0}(-21,1034)(5,1034)(5,1047)(-10,1047)(-10,1032)(0,1032){1}
wire w166;    //: /sn:0 {0}(5,532)(-17,532)(-17,676){1}
wire w134;    //: /sn:0 {0}(-3020,359)(-3020,79)(-3019,79)(-3019,71){1}
wire w122;    //: /sn:0 {0}(-2584,399)(-2584,1289)(-276,1289)(-276,1321){1}
wire w244;    //: /sn:0 {0}(-257,1379)(-257,1486)(-239,1486)(-239,1501){1}
wire w220;    //: /sn:0 {0}(-45,1216)(-45,1305)(-41,1305)(-41,1320){1}
wire w141;    //: /sn:0 {0}(377,556)(377,664)(383,664)(383,679){1}
wire w14;    //: /sn:0 {0}(364,397)(364,483)(309,483)(309,498){1}
wire w56;    //: /sn:0 {0}(-774,354)(-774,320)(-721,320){1}
//: {2}(-717,320)(-665,320){3}
//: {4}(-661,320)(-608,320){5}
//: {6}(-604,320)(-552,320){7}
//: {8}(-548,320)(-501,320){9}
//: {10}(-497,320)(-446,320){11}
//: {12}(-442,320)(-392,320){13}
//: {14}(-390,318)(-390,108)(-392,108)(-392,102){15}
//: {16}(-390,322)(-390,355){17}
//: {18}(-444,322)(-444,334)(-443,334)(-443,355){19}
//: {20}(-499,322)(-499,332)(-498,332)(-498,355){21}
//: {22}(-550,322)(-550,332)(-551,332)(-551,354){23}
//: {24}(-606,322)(-606,354){25}
//: {26}(-663,322)(-663,354){27}
//: {28}(-719,322)(-719,354){29}
wire w16;    //: /sn:0 {0}(-410,355)(-410,79)(-413,79)(-413,71){1}
wire w179;    //: /sn:0 {0}(-4,710)(14,710)(14,706)(16,706){1}
wire w81;    //: /sn:0 {0}(-1864,357)(-1864,79)(-1866,79)(-1866,71){1}
wire w89;    //: /sn:0 {0}(-1721,356)(-1721,71){1}
wire w19;    //: /sn:0 {0}(9,397)(9,420)(430,420)(430,498){1}
wire w4;    //: /sn:0 {0}(51,355)(51,79)(50,79)(50,71){1}
wire w195;    //: /sn:0 {0}(-91,891)(-73,891)(-73,888)(-68,888){1}
wire w38;    //: /sn:0 {0}(-324,355)(-324,213)(-326,213)(-326,71){1}
wire w182;    //: /sn:0 {0}(160,917)(160,985)(166,985)(166,1000){1}
wire w180;    //: /sn:0 {0}(42,734)(42,843)(33,843)(33,858){1}
wire w152;    //: /sn:0 {0}(301,556)(301,664)(317,664)(317,679){1}
wire w183;    //: /sn:0 {0}(-51,706)(-104,706)(-104,857){1}
wire w194;    //: /sn:0 {0}(162,1216)(162,1321){1}
wire w181;    //: /sn:0 {0}(-783,396)(-783,670)(-44,670)(-44,676){1}
wire w3;    //: /sn:0 {0}(516,355)(516,71){1}
wire w0;    //: /sn:0 {0}(569,355)(569,71){1}
wire w151;    //: /sn:0 {0}(253,532)(267,532)(267,528)(275,528){1}
wire w128;    //: /sn:0 {0}(-2912,359)(-2912,79)(-2913,79)(-2913,71){1}
wire w127;    //: /sn:0 {0}(-2847,400)(-2847,1407)(-69,1407)(-69,1501){1}
wire w120;    //: /sn:0 {0}(-2595,357)(-2595,79)(-2594,79)(-2594,71){1}
wire w240;    //: /sn:0 {0}(-189,1380)(-189,1486)(-174,1486)(-174,1501){1}
wire w133;    //: /sn:0 {0}(-2956,401)(-2956,1428)(-201,1428)(-201,1501){1}
wire w111;    //: /sn:0 {0}(-2439,357)(-2439,79)(-2438,79)(-2438,71){1}
wire w104;    //: /sn:0 {0}(-2324,399)(-2324,1237)(72,1237)(72,1320){1}
wire w168;    //: /sn:0 {0}(242,736)(242,844)(235,844)(235,859){1}
wire w171;    //: /sn:0 {0}(128,710)(139,710)(139,707)(139,707)(139,707)(149,707){1}
wire w204;    //: /sn:0 {0}(26,1060)(26,1143)(31,1143)(31,1158){1}
wire w75;    //: /sn:0 {0}(-2115,357)(-2115,335)(-2113,335)(-2113,325){1}
//: {2}(-2111,323)(-2063,323){3}
//: {4}(-2059,323)(-2007,323){5}
//: {6}(-2003,323)(-1953,323){7}
//: {8}(-1949,323)(-1900,323){9}
//: {10}(-1896,323)(-1844,323){11}
//: {12}(-1840,323)(-1794,323){13}
//: {14}(-1792,321)(-1792,108)(-1793,108)(-1793,102){15}
//: {16}(-1792,325)(-1792,357){17}
//: {18}(-1842,325)(-1842,346)(-1844,346)(-1844,357){19}
//: {20}(-1898,325)(-1898,335)(-1897,335)(-1897,357){21}
//: {22}(-1951,325)(-1951,335)(-1952,335)(-1952,357){23}
//: {24}(-2005,325)(-2005,357){25}
//: {26}(-2061,325)(-2061,357){27}
//: {28}(-2115,323)(-2168,323)(-2168,357){29}
wire w237;    //: /sn:0 {0}(-95,1535)(-71,1535)(-71,1531)(-76,1531){1}
wire w209;    //: /sn:0 {0}(42,1354)(58,1354)(58,1350)(65,1350){1}
wire w119;    //: /sn:0 {0}(-2533,399)(-2533,1279)(-208,1279)(-208,1322){1}
wire w67;    //: /sn:0 {0}(-1812,357)(-1812,79)(-1813,79)(-1813,71){1}
wire w54;    //: /sn:0 {0}(-728,396)(-728,663)(23,663)(23,676){1}
wire w215;    //: /sn:0 {0}(-201,1030)(-242,1030)(-242,1157){1}
wire w90;    //: /sn:0 {0}(-1917,357)(-1917,79)(-1918,79)(-1918,71){1}
wire w176;    //: /sn:0 {0}(107,734)(107,844)(99,844)(99,859){1}
wire w156;    //: /sn:0 {0}(232,556)(232,663)(250,663)(250,678){1}
wire w167;    //: /sn:0 {0}(27,555)(27,661)(50,661)(50,676){1}
wire w36;    //: /sn:0 {0}(-452,397)(-452,624)(356,624)(356,679){1}
wire w41;    //: /sn:0 {0}(-1184,356)(-1184,325){1}
//: {2}(-1182,323)(-1131,323){3}
//: {4}(-1127,323)(-1075,323){5}
//: {6}(-1071,323)(-1022,323){7}
//: {8}(-1018,323)(-968,323){9}
//: {10}(-964,323)(-912,323){11}
//: {12}(-908,323)(-857,323){13}
//: {14}(-855,321)(-855,108)(-857,108)(-857,102){15}
//: {16}(-855,325)(-855,355){17}
//: {18}(-910,325)(-910,355){19}
//: {20}(-966,325)(-966,335)(-965,335)(-965,355){21}
//: {22}(-1020,325)(-1020,335)(-1019,335)(-1019,355){23}
//: {24}(-1073,325)(-1073,335)(-1074,335)(-1074,355){25}
//: {26}(-1129,325)(-1129,356){27}
//: {28}(-1186,323)(-1238,323)(-1238,356){29}
wire w124;    //: /sn:0 {0}(-2858,358)(-2858,79)(-2859,79)(-2859,71){1}
wire w23;    //: /sn:0 {0}(200,396)(200,475)(100,475)(100,498){1}
wire w20;    //: /sn:0 {0}(255,396)(255,479)(169,479)(169,498){1}
wire w174;    //: /sn:0 {0}(179,1034)(200,1034)(200,1030)(200,1030){1}
wire w108;    //: /sn:0 {0}(-2177,399)(-2177,1125)(-269,1125)(-269,1157){1}
wire w225;    //: /sn:0 {0}(-29,1535)(14,1535)(14,1530)(-5,1530){1}
wire w82;    //: /sn:0 {0}(-1549,398)(-1549,959)(7,959)(7,1002){1}
wire w126;    //: /sn:0 {0}(-399,397)(-399,615)(429,615)(429,680){1}
wire w223;    //: /sn:0 {0}(-162,1191)(-145,1191)(-145,1188)(-141,1188){1}
wire w158;    //: /sn:0 {0}(309,737)(309,844)(307,844)(307,859){1}
wire w74;    //: /sn:0 {0}(-1247,398)(-1247,852)(-131,852)(-131,857){1}
wire w125;    //: /sn:0 {0}(-2636,399)(-2636,1306)(-341,1306)(-341,1321){1}
wire w35;    //: /sn:0 {0}(-270,355)(-270,71){1}
wire w91;    //: /sn:0 {0}(-1710,398)(-1710,985)(-194,985)(-194,1000){1}
wire w103;    //: /sn:0 {0}(-2135,357)(-2135,79)(-2136,79)(-2136,71){1}
wire w8;    //: /sn:0 {0}(472,397)(472,483)(457,483)(457,498){1}
wire w192;    //: /sn:0 {0}(25,916)(25,987)(34,987)(34,1002){1}
wire w163;    //: /sn:0 {0}(35,499)(35,486)(66,486)(66,528)(66,528){1}
wire w101;    //: /sn:0 {0}(-2748,358)(-2748,79)(-2751,79)(-2751,71){1}
wire w71;    //: /sn:0 {0}(-1193,398)(-1193,846)(-61,846)(-61,858){1}
wire w238;    //: /sn:0 {0}(63,1797)(63,1602)(-50,1602)(-50,1559){1}
wire w144;    //: /sn:0 {0}(449,556)(449,665)(448,665)(448,680){1}
wire w22;    //: /sn:0 {0}(-57,355)(-57,79)(-59,79)(-59,71){1}
wire w17;    //: /sn:0 {0}(310,397)(310,483)(240,483)(240,498){1}
wire w117;    //: /sn:0 {0}(-2544,357)(-2544,79)(-2547,79)(-2547,71){1}
wire w84;    //: /sn:0 {0}(-2284,357)(-2284,71){1}
wire w53;    //: /sn:0 {0}(-919,397)(-919,809)(280,809)(280,859){1}
wire w172;    //: /sn:0 {0}(175,735)(175,844)(168,844)(168,859){1}
wire w263;    //: /sn:0 {0}(3,1797)(3,1666)(-427,1666)(-427,1531)(-411,1531){1}
wire w255;    //: /sn:0 {0}(-294,1535)(-273,1535)(-273,1531)(-273,1531){1}
wire w211;    //: /sn:0 {0}(-154,1034)(-139,1034)(-139,1030)(-135,1030){1}
wire w228;    //: /sn:0 {0}(-183,1215)(-183,1307)(-181,1307)(-181,1322){1}
wire w12;    //: /sn:0 {0}(353,355)(353,79)(352,79)(352,71){1}
wire w113;    //: /sn:0 {0}(-2428,399)(-2428,1256)(-68,1256)(-68,1320){1}
wire w44;    //: /sn:0 {0}(-864,397)(-864,801)(357,801)(357,860){1}
wire w2;    //: /sn:0 {0}(580,397)(580,1782)(153,1782)(153,1797){1}
wire w226;    //: /sn:0 {0}(73,1797)(73,1573)(21,1573)(21,1558){1}
wire w115;    //: /sn:0 {0}(-2804,358)(-2804,79)(-2805,79)(-2805,71){1}
wire w83;    //: /sn:0 {0}(-1614,356)(-1614,79)(-1615,79)(-1615,71){1}
wire w77;    //: /sn:0 {0}(-1506,356)(-1506,79)(-1505,79)(-1505,71){1}
wire w200;    //: /sn:0 {0}(-112,915)(-112,985)(-101,985)(-101,1000){1}
wire w78;    //: /sn:0 {0}(-1801,399)(-1801,1068)(215,1068)(215,1159){1}
wire w10;    //: /sn:0 {0}(62,397)(62,410)(506,410)(506,499){1}
wire w224;    //: /sn:0 {0}(-115,1216)(-115,1306)(-111,1306)(-111,1321){1}
wire w190;    //: /sn:0 {0}(158,1058)(158,1143)(170,1143)(170,1158){1}
wire w246;    //: /sn:0 {0}(53,1797)(53,1611)(-116,1611)(-116,1559){1}
wire w138;    //: /sn:0 {0}(440,736)(440,1769)(133,1769)(133,1797){1}
wire w86;    //: /sn:0 {0}(-1668,356)(-1668,79)(-1667,79)(-1667,71){1}
wire w95;    //: /sn:0 {0}(-2273,399)(-2273,1230)(143,1230)(143,1321){1}
wire w52;    //: /sn:0 {0}(-739,354)(-739,71){1}
wire w188;    //: /sn:0 {0}(91,917)(91,985)(99,985)(99,1000){1}
wire w231;    //: /sn:0 {0}(-276,1187)(-314,1187)(-314,1321){1}
wire w29;    //: /sn:0 {0}(-163,355)(-163,79)(-164,79)(-164,71){1}
wire w80;    //: /sn:0 {0}(-1560,356)(-1560,79)(-1561,79)(-1561,71){1}
wire w142;    //: /sn:0 {0}(-3116,400)(-3116,1486)(-404,1486)(-404,1501){1}
wire w155;    //: /sn:0 {0}(182,532)(204,532)(204,528)(206,528){1}
wire w178;    //: /sn:0 {0}(112,893)(127,893)(127,889)(134,889){1}
wire w187;    //: /sn:0 {0}(46,892)(62,892)(62,889)(65,889){1}
wire w147;    //: /sn:0 {0}(322,532)(336,532)(336,528)(351,528){1}
wire w42;    //: /sn:0 {0}(-507,397)(-507,633)(290,633)(290,679){1}
wire w264;    //: /sn:0 {0}(13,1797)(13,1652)(-385,1652)(-385,1559){1}
wire w50;    //: /sn:0 {0}(-1344,356)(-1344,79)(-1343,79)(-1343,71){1}
wire w6;    //: /sn:0 {0}(461,355)(461,71){1}
wire w247;    //: /sn:0 {0}(-348,1351)(-377,1351)(-377,1501){1}
wire w93;    //: /sn:0 {0}(-1906,399)(-1906,1083)(76,1083)(76,1158){1}
wire w7;    //: /sn:0 {0}(-250,355)(-250,336)(-251,336)(-251,326){1}
//: {2}(-249,324)(-198,324){3}
//: {4}(-194,324)(-144,324){5}
//: {6}(-140,324)(-92,324){7}
//: {8}(-88,324)(-38,324){9}
//: {10}(-34,324)(16,324){11}
//: {12}(20,324)(69,324){13}
//: {14}(71,322)(71,108)(70,108)(70,102){15}
//: {16}(71,326)(71,355){17}
//: {18}(18,326)(18,355){19}
//: {20}(-36,326)(-36,336)(-37,336)(-37,355){21}
//: {22}(-90,326)(-90,355){23}
//: {24}(-142,326)(-142,336)(-143,336)(-143,355){25}
//: {26}(-196,326)(-196,355){27}
//: {28}(-253,324)(-304,324)(-304,355){29}
wire w60;    //: /sn:0 {0}(-1039,355)(-1039,79)(-1042,79)(-1042,71){1}
wire w112;    //: /sn:0 {0}(-2737,400)(-2737,1391)(74,1391)(74,1500){1}
wire w99;    //: /sn:0 {0}(-2014,399)(-2014,1097)(-64,1097)(-64,1158){1}
wire w61;    //: /sn:0 {0}(-1333,398)(-1333,927)(279,927)(279,1001){1}
wire w175;    //: /sn:0 {0}(63,710)(81,710)(81,706)(81,706){1}
wire w46;    //: /sn:0 {0}(-626,354)(-626,71){1}
wire w135;    //: /sn:0 {0}(396,713)(413,713)(413,713)(418,713){1}
wire w153;    //: /sn:0 {0}(248,893)(281,893)(281,889)(273,889){1}
wire w15;    //: /sn:0 {0}(299,355)(299,79)(297,79)(297,71){1}
wire w216;    //: /sn:0 {0}(-175,1058)(-175,1157){1}
wire w129;    //: /sn:0 {0}(470,532)(497,532)(497,532)(495,532){1}
wire w109;    //: /sn:0 {0}(-3053,359)(-3053,327){1}
//: {2}(-3051,325)(-3003,325){3}
//: {4}(-2999,325)(-2949,325){5}
//: {6}(-2945,325)(-2894,325){7}
//: {8}(-2890,325)(-2841,325){9}
//: {10}(-2837,325)(-2787,325){11}
//: {12}(-2783,325)(-2730,325){13}
//: {14}(-2728,323)(-2728,102){15}
//: {16}(-2728,327)(-2728,358){17}
//: {18}(-2785,327)(-2785,347)(-2784,347)(-2784,358){19}
//: {20}(-2839,327)(-2839,337)(-2838,337)(-2838,358){21}
//: {22}(-2892,327)(-2892,359){23}
//: {24}(-2947,327)(-2947,359){25}
//: {26}(-3001,327)(-3001,337)(-3000,337)(-3000,359){27}
//: {28}(-3055,325)(-3107,325)(-3107,358){29}
wire w106;    //: /sn:0 {0}(-2188,357)(-2188,71){1}
wire w69;    //: /sn:0 {0}(-1204,356)(-1204,71){1}
wire w51;    //: /sn:0 {0}(-672,396)(-672,655)(88,655)(88,676){1}
wire w207;    //: /sn:0 {0}(-88,1034)(-68,1034)(-68,1030)(-68,1030){1}
wire w213;    //: /sn:0 {0}(-24,1192)(-11,1192)(-11,1188)(-3,1188){1}
wire w239;    //: /sn:0 {0}(-236,1355)(-224,1355)(-224,1352)(-215,1352){1}
wire w229;    //: /sn:0 {0}(-98,1355)(-79,1355)(-79,1350)(-75,1350){1}
wire w97;    //: /sn:0 {0}(-2025,357)(-2025,79)(-2026,79)(-2026,71){1}
wire w114;    //: /sn:0 {0}(-2492,357)(-2492,71){1}
wire w245;    //: /sn:0 {0}(-161,1535)(-148,1535)(-148,1531)(-142,1531){1}
wire w64;    //: /sn:0 {0}(-1397,356)(-1397,79)(-1401,79)(-1401,71){1}
wire w66;    //: /sn:0 {0}(-1149,356)(-1149,79)(-1150,79)(-1150,71){1}
wire w37;    //: /sn:0 {0}(-259,397)(-259,457)(73,457)(73,498){1}
wire w177;    //: /sn:0 {0}(226,1058)(226,1144)(234,1144)(234,1159){1}
wire w159;    //: /sn:0 {0}(113,532)(137,532)(137,528)(135,528){1}
wire w63;    //: /sn:0 {0}(-1094,355)(-1094,71){1}
wire w259;    //: /sn:0 {0}(-364,1535)(-353,1535)(-353,1531)(-341,1531){1}
wire w34;    //: /sn:0 {0}(-205,397)(-205,450)(142,450)(142,498){1}
wire w236;    //: /sn:0 {0}(-119,1379)(-119,1486)(-108,1486)(-108,1501){1}
wire w21;    //: /sn:0 {0}(189,354)(189,79)(187,79)(187,71){1}
wire w76;    //: /sn:0 {0}(-1440,398)(-1440,942)(139,942)(139,1000){1}
wire w102;    //: /sn:0 {0}(-2070,399)(-2070,1105)(-134,1105)(-134,1158){1}
wire w87;    //: /sn:0 {0}(-1853,399)(-1853,1075)(143,1075)(143,1158){1}
wire w43;    //: /sn:0 {0}(-571,354)(-571,79)(-574,79)(-574,71){1}
wire w157;    //: /sn:0 {0}(263,712)(294,712)(294,709)(283,709){1}
wire w199;    //: /sn:0 {0}(-138,887)(-167,887)(-167,1000){1}
wire w170;    //: /sn:0 {0}(92,556)(92,661)(115,661)(115,676){1}
wire w230;    //: /sn:0 {0}(-49,1378)(-49,1486)(-42,1486)(-42,1501){1}
wire w31;    //: /sn:0 {0}(-152,397)(-152,444)(213,444)(213,498){1}
wire w100;    //: /sn:0 {0}(-2081,357)(-2081,79)(-2080,79)(-2080,71){1}
wire w58;    //: /sn:0 {0}(-1648,356)(-1648,335)(-1649,335)(-1649,325){1}
//: {2}(-1647,323)(-1595,323){3}
//: {4}(-1591,323)(-1541,323){5}
//: {6}(-1537,323)(-1488,323){7}
//: {8}(-1484,323)(-1432,323){9}
//: {10}(-1428,323)(-1379,323){11}
//: {12}(-1375,323)(-1326,323){13}
//: {14}(-1324,321)(-1324,102){15}
//: {16}(-1324,325)(-1324,356){17}
//: {18}(-1377,325)(-1377,356){19}
//: {20}(-1430,325)(-1430,335)(-1431,335)(-1431,356){21}
//: {22}(-1486,325)(-1486,356){23}
//: {24}(-1539,325)(-1539,335)(-1540,335)(-1540,356){25}
//: {26}(-1593,325)(-1593,335)(-1594,335)(-1594,356){27}
//: {28}(-1651,323)(-1701,323)(-1701,356){29}
wire w130;    //: /sn:0 {0}(-2901,401)(-2901,1418)(-135,1418)(-135,1501){1}
wire w169;    //: /sn:0 {0}(-615,396)(-615,648)(156,648)(156,677){1}
wire w28;    //: /sn:0 {0}(-99,397)(-99,437)(282,437)(282,498){1}
wire w251;    //: /sn:0 {0}(-226,1535)(-210,1535)(-210,1531)(-208,1531){1}
wire w24;    //: /sn:0 {0}(-793,71)(-793,79)(-794,79)(-794,354){1}
wire w161;    //: /sn:0 {0}(226,1215)(226,1742)(103,1742)(103,1797){1}
wire w1;    //: /sn:0 {0}(264,354)(264,329)(263,329)(263,319){1}
//: {2}(265,317)(315,317){3}
//: {4}(319,317)(370,317){5}
//: {6}(374,317)(424,317){7}
//: {8}(428,317)(477,317){9}
//: {10}(481,317)(533,317){11}
//: {12}(537,317)(587,317){13}
//: {14}(589,315)(589,102){15}
//: {16}(589,319)(589,355){17}
//: {18}(535,319)(535,329)(536,329)(536,355){19}
//: {20}(479,319)(479,329)(481,329)(481,355){21}
//: {22}(426,319)(426,329)(428,329)(428,355){23}
//: {24}(372,319)(372,329)(373,329)(373,355){25}
//: {26}(317,319)(317,329)(319,329)(319,355){27}
//: {28}(261,317)(209,317)(209,354){29}
wire w256;    //: /sn:0 {0}(33,1797)(33,1630)(-247,1630)(-247,1559){1}
wire w260;    //: /sn:0 {0}(23,1797)(23,1640)(-315,1640)(-315,1559){1}
wire w184;    //: /sn:0 {0}(-25,734)(-25,843)(-34,843)(-34,858){1}
wire w132;    //: /sn:0 {0}(517,555)(517,1774)(143,1774)(143,1797){1}
wire w235;    //: /sn:0 {0}(-168,1356)(-155,1356)(-155,1351)(-145,1351){1}
wire w221;    //: /sn:0 {0}(-28,1354)(-10,1354)(-10,1350)(-5,1350){1}
wire w196;    //: /sn:0 {0}(-42,916)(-42,985)(-34,985)(-34,1000){1}
wire w140;    //: /sn:0 {0}(-3127,358)(-3127,79)(-3128,79)(-3128,71){1}
wire w205;    //: /sn:0 {0}(44,1192)(65,1192)(65,1188)(69,1188){1}
wire w154;    //: /sn:0 {0}(299,917)(299,986)(298,986)(298,1001){1}
wire w25;    //: /sn:0 {0}(-46,397)(-46,429)(358,429)(358,498){1}
wire w227;    //: /sn:0 {0}(-229,1191)(-213,1191)(-213,1187)(-209,1187){1}
wire w116;    //: /sn:0 {0}(-2481,399)(-2481,1270)(-138,1270)(-138,1321){1}
wire w98;    //: /sn:0 {0}(-2335,357)(-2335,71){1}
wire w65;    //: /sn:0 {0}(-1083,397)(-1083,832)(72,832)(72,859){1}
wire w210;    //: /sn:0 {0}(91,1378)(91,1485)(93,1485)(93,1500){1}
wire w243;    //: /sn:0 {0}(-301,1355)(-283,1355)(-283,1351)(-283,1351){1}
wire w212;    //: /sn:0 {0}(-109,1058)(-109,1143)(-107,1143)(-107,1158){1}
wire w118;    //: /sn:0 {0}(368,916)(368,1761)(123,1761)(123,1797){1}
wire w18;    //: /sn:0 {0}(244,354)(244,79)(247,79)(247,71){1}
wire w40;    //: /sn:0 {0}(-313,397)(-313,467)(16,467)(16,499){1}
wire w92;    //: /sn:0 {0}(-2575,357)(-2575,327){1}
//: {2}(-2573,325)(-2528,325){3}
//: {4}(-2524,325)(-2474,325){5}
//: {6}(-2470,325)(-2421,325){7}
//: {8}(-2417,325)(-2368,325){9}
//: {10}(-2364,325)(-2316,325){11}
//: {12}(-2312,325)(-2266,325){13}
//: {14}(-2264,323)(-2264,108)(-2265,108)(-2265,102){15}
//: {16}(-2264,327)(-2264,357){17}
//: {18}(-2314,327)(-2314,346)(-2315,346)(-2315,357){19}
//: {20}(-2366,327)(-2366,337)(-2367,337)(-2367,357){21}
//: {22}(-2419,327)(-2419,357){23}
//: {24}(-2472,327)(-2472,357){25}
//: {26}(-2526,327)(-2526,337)(-2524,337)(-2524,357){27}
//: {28}(-2577,325)(-2627,325)(-2627,357){29}
wire w121;    //: /sn:0 {0}(-2793,400)(-2793,1399)(2,1399)(2,1500){1}
wire w164;    //: /sn:0 {0}(181,893)(198,893)(198,889)(201,889){1}
wire w68;    //: /sn:0 {0}(-1138,398)(-1138,838)(6,838)(6,858){1}
wire w30;    //: /sn:0 {0}(-463,355)(-463,79)(-464,79)(-464,71){1}
wire w162;    //: /sn:0 {0}(112,1354)(129,1354)(129,1354)(132,1354){1}
wire w198;    //: /sn:0 {0}(91,1058)(91,1143)(103,1143)(103,1158){1}
wire w149;    //: /sn:0 {0}(330,713)(355,713)(355,709)(349,709){1}
wire w146;    //: /sn:0 {0}(290,1057)(290,1752)(113,1752)(113,1797){1}
wire w222;    //: /sn:0 {0}(21,1378)(21,1485)(29,1485)(29,1500){1}
wire w123;    //: /sn:0 {0}(-2647,357)(-2647,79)(-2649,79)(-2649,71){1}
wire w59;    //: /sn:0 {0}(-974,397)(-974,818)(208,818)(208,859){1}
wire w165;    //: /sn:0 {0}(196,711)(212,711)(212,708)(216,708){1}
wire w185;    //: /sn:0 {0}(154,1377)(154,1734)(93,1734)(93,1797){1}
wire w85;    //: /sn:0 {0}(-1603,398)(-1603,969)(-61,969)(-61,1000){1}
wire w62;    //: /sn:0 {0}(-1028,397)(-1028,826)(141,826)(141,859){1}
wire w248;    //: /sn:0 {0}(-322,1379)(-322,1486)(-307,1486)(-307,1501){1}
wire w197;    //: /sn:0 {0}(47,1036)(55,1036)(55,1030)(55,1030)(55,1030)(65,1030){1}
wire w11;    //: /sn:0 {0}(419,397)(419,483)(385,483)(385,498){1}
wire w137;    //: /sn:0 {0}(-3073,359)(-3073,71){1}
wire w139;    //: /sn:0 {0}(-3062,401)(-3062,1447)(-334,1447)(-334,1501){1}
wire w136;    //: /sn:0 {0}(-3009,401)(-3009,1438)(-266,1438)(-266,1501){1}
wire w49;    //: /sn:0 {0}(-683,354)(-683,79)(-684,79)(-684,71){1}
wire w57;    //: /sn:0 {0}(320,893)(344,893)(344,893)(346,893){1}
wire w173;    //: /sn:0 {0}(227,917)(227,985)(234,985)(234,1000){1}
wire w193;    //: /sn:0 {0}(116,1192)(139,1192)(139,1188)(136,1188){1}
wire w189;    //: /sn:0 {0}(112,1034)(129,1034)(129,1030)(132,1030){1}
wire w110;    //: /sn:0 {0}(-2376,399)(-2376,1245)(2,1245)(2,1320){1}
wire w70;    //: /sn:0 {0}(-1386,398)(-1386,934)(207,934)(207,1000){1}
wire w150;    //: /sn:0 {0}(375,737)(375,845)(376,845)(376,860){1}
wire w105;    //: /sn:0 {0}(-2124,399)(-2124,1113)(-202,1113)(-202,1157){1}
wire w148;    //: /sn:0 {0}(204,1192)(199,1192)(199,1192)(183,1192){1}
wire w252;    //: /sn:0 {0}(43,1797)(43,1620)(-182,1620)(-182,1559){1}
wire w206;    //: /sn:0 {0}(95,1216)(95,1305)(99,1305)(99,1320){1}
wire w186;    //: /sn:0 {0}(42,1534)(58,1534)(58,1533)(63,1533){1}
wire w88;    //: /sn:0 {0}(-1657,398)(-1657,975)(-128,975)(-128,1000){1}
wire w13;    //: /sn:0 {0}(-2,355)(-2,79)(-3,79)(-3,71){1}
wire w72;    //: /sn:0 {0}(-1258,356)(-1258,79)(-1260,79)(-1260,71){1}
wire w94;    //: /sn:0 {0}(-1972,357)(-1972,79)(-1974,79)(-1974,71){1}
wire w208;    //: /sn:0 {0}(-42,1058)(-42,1143)(-37,1143)(-37,1158){1}
wire w5;    //: /sn:0 {0}(527,397)(527,484)(525,484)(525,499){1}
wire w33;    //: /sn:0 {0}(-875,355)(-875,79)(-877,79)(-877,71){1}
wire w191;    //: /sn:0 {0}(-21,892)(4,892)(4,888)(-1,888){1}
wire w47;    //: /sn:0 {0}(-930,355)(-930,79)(-928,79)(-928,71){1}
wire w131;    //: /sn:0 {0}(-2967,359)(-2967,79)(-2969,79)(-2969,71){1}
wire w143;    //: /sn:0 {0}(398,532)(414,532)(414,528)(423,528){1}
wire w107;    //: /sn:0 {0}(-2387,357)(-2387,79)(-2388,79)(-2388,71){1}
wire w9;    //: /sn:0 {0}(408,355)(408,71){1}
wire w79;    //: /sn:0 {0}(-1495,398)(-1495,950)(72,950)(72,1000){1}
wire w145;    //: /sn:0 {0}(247,1034)(275,1034)(275,1034)(268,1034){1}
wire w219;    //: /sn:0 {0}(-94,1192)(-77,1192)(-77,1188)(-71,1188){1}
wire w26;    //: /sn:0 {0}(-110,355)(-110,79)(-112,79)(-112,71){1}
wire w201;    //: /sn:0 {0}(83,1797)(83,1571)(85,1571)(85,1556){1}
wire w232;    //: /sn:0 {0}(-250,1215)(-250,1306)(-249,1306)(-249,1321){1}
wire w39;    //: /sn:0 {0}(-518,355)(-518,79)(-519,79)(-519,71){1}
wire w55;    //: /sn:0 {0}(-985,355)(-985,79)(-986,79)(-986,71){1}
//: enddecls

  FA g237 (.B(w220), .A(w113), .Cin(w221), .Cout(w229), .S(w230));   //: @(-74, 1321) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w111 = A[3]; //: TAP g165 @(-2438,65) /sn:0 /R:1 /w:[ 1 104 103 ] /ss:1
  AND2 g154 (.in1(w92), .in2(w123), .out(w125));   //: @(-2657, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  AND2 g4 (.in1(w1), .in2(w6), .out(w8));   //: @(451, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  AND2 g8 (.in1(w1), .in2(w18), .out(w20));   //: @(234, 355) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  assign w101 = A[0]; //: TAP g186 @(-2751,65) /sn:0 /R:1 /w:[ 1 114 113 ] /ss:1
  assign w90 = A[2]; //: TAP g140 @(-1918,65) /sn:0 /R:1 /w:[ 1 86 85 ] /ss:1
  //: joint g13 (w1) @(479, 317) /w:[ 10 -1 9 20 ]
  //: joint g37 (w7) @(18, 324) /w:[ 12 -1 11 18 ]
  AND2 g55 (.in1(w56), .in2(w49), .out(w51));   //: @(-693, 355) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  assign w56 = B[2]; //: TAP g58 @(-392,96) /sn:0 /R:1 /w:[ 15 6 5 ] /ss:1
  assign w81 = A[1]; //: TAP g139 @(-1866,65) /sn:0 /R:1 /w:[ 1 84 83 ] /ss:1
  //: joint g112 (w58) @(-1593, 323) /w:[ 4 -1 3 26 ]
  FA g211 (.B(w158), .A(w53), .Cin(w57), .Cout(w153), .S(w154));   //: @(274, 860) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  AND2 g76 (.in1(w41), .in2(w55), .out(w59));   //: @(-995, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  //: joint g111 (w58) @(-1539, 323) /w:[ 6 -1 5 24 ]
  HA g218 (.B(w154), .A(w61), .Cout(w145), .S(w146));   //: @(269, 1002) /sz:(40, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  AND2 g176 (.in1(w109), .in2(w137), .out(w139));   //: @(-3083, 360) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  //: joint g157 (w92) @(-2366, 325) /w:[ 10 -1 9 20 ]
  FA g238 (.B(w224), .A(w116), .Cin(w229), .Cout(w235), .S(w236));   //: @(-144, 1322) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w98 = A[1]; //: TAP g163 @(-2335,65) /sn:0 /R:1 /w:[ 1 100 99 ] /ss:1
  //: IN g1 (B) @(617,98) /sn:0 /R:2 /w:[ 0 ]
  //: joint g64 (w56) @(-663, 320) /w:[ 4 -1 3 26 ]
  assign w114 = A[4]; //: TAP g166 @(-2492,65) /sn:0 /R:1 /w:[ 1 106 105 ] /ss:1
  //: joint g11 (w1) @(589, 317) /w:[ -1 14 13 16 ]
  FA g241 (.B(w231), .A(w125), .Cin(w243), .Cout(w247), .S(w248));   //: @(-347, 1322) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  FA g206 (.A(w169), .B(w160), .Cin(w165), .Cout(w171), .S(w172));   //: @(150, 678) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  AND2 g130 (.in1(w75), .in2(w106), .out(w108));   //: @(-2198, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  assign w89 = A[7]; //: TAP g121 @(-1721,65) /sn:0 /R:1 /w:[ 1 80 79 ] /ss:1
  AND2 g28 (.in1(w7), .in2(w22), .out(w25));   //: @(-67, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  AND2 g50 (.in1(w56), .in2(w16), .out(w126));   //: @(-420, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  FA g223 (.B(w196), .A(w85), .Cin(w203), .Cout(w207), .S(w208));   //: @(-67, 1001) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g197 (.A(w28), .B(w14), .Cin(w147), .Cout(w151), .S(w152));   //: @(276, 499) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g132 (w75) @(-1842, 323) /w:[ 12 -1 11 18 ]
  assign w3 = A[1]; //: TAP g19 @(516,65) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: joint g113 (w58) @(-1649, 323) /w:[ 2 -1 28 1 ]
  FA g225 (.B(w199), .A(w91), .Cin(w211), .Cout(w215), .S(w216));   //: @(-200, 1001) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  AND2 g150 (.in1(w92), .in2(w111), .out(w113));   //: @(-2449, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  AND2 g146 (.in1(w92), .in2(w84), .out(w95));   //: @(-2294, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  FA g208 (.A(w54), .B(w167), .Cin(w175), .Cout(w179), .S(w180));   //: @(17, 677) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w137 = A[6]; //: TAP g192 @(-3073,65) /sn:0 /R:1 /w:[ 1 126 125 ] /ss:1
  AND2 g177 (.in1(w109), .in2(w140), .out(w142));   //: @(-3137, 359) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  AND2 g6 (.in1(w1), .in2(w12), .out(w14));   //: @(343, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  //: joint g38 (w7) @(-36, 324) /w:[ 10 -1 9 20 ]
  assign w64 = A[1]; //: TAP g115 @(-1401,65) /sn:0 /R:1 /w:[ 1 68 67 ] /ss:1
  AND2 g7 (.in1(w1), .in2(w15), .out(w17));   //: @(289, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  AND2 g53 (.in1(w56), .in2(w43), .out(w45));   //: @(-581, 355) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  AND2 g75 (.in1(w41), .in2(w47), .out(w53));   //: @(-940, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  FA g227 (.B(w190), .A(w87), .Cin(w148), .Cout(w193), .S(w194));   //: @(137, 1159) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  assign w123 = A[7]; //: TAP g169 @(-2649,65) /sn:0 /R:1 /w:[ 1 112 111 ] /ss:1
  //: joint g160 (w92) @(-2526, 325) /w:[ 4 -1 3 26 ]
  //: joint g135 (w75) @(-2005, 323) /w:[ 6 -1 5 24 ]
  assign w6 = A[2]; //: TAP g20 @(461,65) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  AND2 g31 (.in1(w7), .in2(w32), .out(w34));   //: @(-226, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  FA g230 (.B(w208), .A(w99), .Cin(w213), .Cout(w219), .S(w220));   //: @(-70, 1159) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  AND2 g149 (.in1(w92), .in2(w107), .out(w110));   //: @(-2397, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  AND2 g124 (.in1(w75), .in2(w90), .out(w93));   //: @(-1927, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  FA g207 (.A(w51), .B(w170), .Cin(w171), .Cout(w175), .S(w176));   //: @(82, 677) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g39 (w7) @(-90, 324) /w:[ 8 -1 7 22 ]
  assign w39 = A[2]; //: TAP g68 @(-519,65) /sn:0 /R:1 /w:[ 1 38 37 ] /ss:1
  FA g200 (.A(w37), .B(w23), .Cin(w159), .Cout(w163), .S(w170));   //: @(67, 499) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w35 = A[6]; //: TAP g48 @(-270,65) /sn:0 /R:1 /w:[ 1 30 29 ] /ss:1
  FA g195 (.A(w19), .B(w8), .Cin(w129), .Cout(w143), .S(w144));   //: @(424, 499) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g17 (w1) @(263, 317) /w:[ 2 -1 28 1 ]
  assign w21 = A[7]; //: TAP g25 @(187,65) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  AND2 g29 (.in1(w7), .in2(w26), .out(w28));   //: @(-120, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  FA g205 (.A(w45), .B(w156), .Cin(w157), .Cout(w165), .S(w168));   //: @(217, 679) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g179 (w109) @(-2728, 325) /w:[ -1 14 13 16 ]
  AND2 g52 (.in1(w56), .in2(w39), .out(w42));   //: @(-528, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  assign w58 = B[4]; //: TAP g106 @(-1324,96) /sn:0 /R:1 /w:[ 15 10 9 ] /ss:1
  //: joint g107 (w58) @(-1324, 323) /w:[ -1 14 13 16 ]
  FA g231 (.B(w212), .A(w102), .Cin(w219), .Cout(w223), .S(w224));   //: @(-140, 1159) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  AND2 g174 (.in1(w109), .in2(w131), .out(w133));   //: @(-2977, 360) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  //: joint g83 (w41) @(-855, 323) /w:[ -1 14 13 16 ]
  FA g221 (.B(w188), .A(w79), .Cin(w189), .Cout(w197), .S(w198));   //: @(66, 1001) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  HA g201 (.A(w40), .B(w163), .Cout(w166), .S(w167));   //: @(6, 500) /sz:(40, 54) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  AND2 g100 (.in1(w58), .in2(w73), .out(w76));   //: @(-1461, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  //: joint g14 (w1) @(426, 317) /w:[ 8 -1 7 22 ]
  FA g248 (.B(w248), .A(w139), .Cin(w255), .Cout(w259), .S(w260));   //: @(-340, 1502) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  HA g202 (.A(w126), .B(w144), .Cout(w135), .S(w138));   //: @(419, 681) /sz:(40, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  assign w140 = A[7]; //: TAP g193 @(-3128,65) /sn:0 /R:1 /w:[ 1 128 127 ] /ss:1
  assign w22 = A[2]; //: TAP g44 @(-59,65) /sn:0 /R:1 /w:[ 1 22 21 ] /ss:1
  assign w32 = A[5]; //: TAP g47 @(-217,65) /sn:0 /R:1 /w:[ 1 28 27 ] /ss:1
  AND2 g80 (.in1(w41), .in2(w69), .out(w71));   //: @(-1214, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  assign w63 = A[4]; //: TAP g94 @(-1094,65) /sn:0 /R:1 /w:[ 1 58 57 ] /ss:1
  FA g247 (.B(w244), .A(w136), .Cin(w251), .Cout(w255), .S(w256));   //: @(-272, 1502) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  FA g232 (.B(w216), .A(w105), .Cin(w223), .Cout(w227), .S(w228));   //: @(-208, 1158) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  AND2 g172 (.in1(w109), .in2(w124), .out(w127));   //: @(-2868, 359) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  //: joint g159 (w92) @(-2472, 325) /w:[ 6 -1 5 24 ]
  assign w9 = A[3]; //: TAP g21 @(408,65) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: joint g84 (w41) @(-910, 323) /w:[ 12 -1 11 18 ]
  AND2 g105 (.in1(w58), .in2(w89), .out(w91));   //: @(-1731, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  FA g236 (.B(w214), .A(w110), .Cin(w209), .Cout(w221), .S(w222));   //: @(-4, 1321) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g155 (w92) @(-2264, 325) /w:[ -1 14 13 16 ]
  assign w94 = A[3]; //: TAP g141 @(-1974,65) /sn:0 /R:1 /w:[ 1 88 87 ] /ss:1
  assign w15 = A[5]; //: TAP g23 @(297,65) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  //: joint g41 (w7) @(-196, 324) /w:[ 4 -1 3 26 ]
  FA g249 (.B(w247), .A(w142), .Cin(w259), .Cout(w263), .S(w264));   //: @(-410, 1502) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  AND2 g151 (.in1(w92), .in2(w114), .out(w116));   //: @(-2502, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  //: joint g40 (w7) @(-142, 324) /w:[ 6 -1 5 24 ]
  AND2 g54 (.in1(w56), .in2(w46), .out(w169));   //: @(-636, 355) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  assign w60 = A[3]; //: TAP g93 @(-1042,65) /sn:0 /R:1 /w:[ 1 56 55 ] /ss:1
  assign w73 = A[2]; //: TAP g116 @(-1453,65) /sn:0 /R:1 /w:[ 1 70 69 ] /ss:1
  AND2 g123 (.in1(w75), .in2(w81), .out(w87));   //: @(-1874, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  FA g222 (.B(w192), .A(w82), .Cin(w197), .Cout(w203), .S(w204));   //: @(1, 1003) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w117 = A[5]; //: TAP g167 @(-2547,65) /sn:0 /R:1 /w:[ 1 108 107 ] /ss:1
  //: IN g0 (A) @(615,67) /sn:0 /R:2 /w:[ 0 ]
  AND2 g26 (.in1(w7), .in2(w4), .out(w10));   //: @(41, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  assign w29 = A[4]; //: TAP g46 @(-164,65) /sn:0 /R:1 /w:[ 1 26 25 ] /ss:1
  assign w33 = A[0]; //: TAP g90 @(-877,65) /sn:0 /R:1 /w:[ 1 50 49 ] /ss:1
  FA g228 (.B(w198), .A(w93), .Cin(w193), .Cout(w205), .S(w206));   //: @(70, 1159) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w41 = B[3]; //: TAP g82 @(-857,96) /sn:0 /R:1 /w:[ 15 8 7 ] /ss:1
  FA g243 (.B(w222), .A(w121), .Cin(w186), .Cout(w225), .S(w226));   //: @(-4, 1501) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  FA g233 (.B(w215), .A(w108), .Cin(w227), .Cout(w231), .S(w232));   //: @(-275, 1158) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  FA g224 (.B(w200), .A(w88), .Cin(w207), .Cout(w211), .S(w212));   //: @(-134, 1001) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g136 (w75) @(-2061, 323) /w:[ 4 -1 3 26 ]
  AND2 g128 (.in1(w75), .in2(w100), .out(w102));   //: @(-2091, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  assign w131 = A[4]; //: TAP g190 @(-2969,65) /sn:0 /R:1 /w:[ 1 122 121 ] /ss:1
  AND2 g173 (.in1(w109), .in2(w128), .out(w130));   //: @(-2922, 360) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  AND2 g33 (.in1(w7), .in2(w38), .out(w40));   //: @(-334, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  assign w47 = A[1]; //: TAP g91 @(-928,65) /sn:0 /R:1 /w:[ 1 52 51 ] /ss:1
  assign w38 = A[7]; //: TAP g49 @(-326,65) /sn:0 /R:1 /w:[ 1 32 31 ] /ss:1
  FA g198 (.A(w31), .B(w17), .Cin(w151), .Cout(w155), .S(w156));   //: @(207, 499) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g137 (w75) @(-2113, 323) /w:[ 2 -1 28 1 ]
  //: joint g61 (w56) @(-499, 320) /w:[ 10 -1 9 20 ]
  AND2 g3 (.in1(w1), .in2(w3), .out(w5));   //: @(506, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  assign w7 = B[1]; //: TAP g34 @(70,96) /sn:0 /R:1 /w:[ 15 4 3 ] /ss:1
  AND2 g51 (.in1(w56), .in2(w30), .out(w36));   //: @(-473, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  //: joint g86 (w41) @(-1020, 323) /w:[ 8 -1 7 22 ]
  //: joint g158 (w92) @(-2419, 325) /w:[ 8 -1 7 22 ]
  FA g220 (.B(w182), .A(w76), .Cin(w174), .Cout(w189), .S(w190));   //: @(133, 1001) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g89 (w41) @(-1184, 323) /w:[ 2 -1 28 1 ]
  FA g217 (.B(w183), .A(w74), .Cin(w195), .Cout(w199), .S(w200));   //: @(-137, 858) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g110 (w58) @(-1486, 323) /w:[ 8 -1 7 22 ]
  AND2 g77 (.in1(w41), .in2(w60), .out(w62));   //: @(-1049, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  //: joint g65 (w56) @(-719, 320) /w:[ 2 -1 1 28 ]
  AND2 g2 (.in1(w1), .in2(w0), .out(w2));   //: @(559, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  assign S = {w263, w264, w260, w256, w252, w246, w238, w226, w201, w185, w161, w146, w118, w138, w132, w2}; //: CONCAT g250  @(78,1802) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g59 (w56) @(-390, 320) /w:[ -1 14 13 16 ]
  assign w92 = B[6]; //: TAP g147 @(-2265,96) /sn:0 /R:1 /w:[ 15 14 13 ] /ss:1
  AND2 g148 (.in1(w92), .in2(w98), .out(w104));   //: @(-2345, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  //: joint g156 (w92) @(-2314, 325) /w:[ 12 -1 11 18 ]
  FA g213 (.B(w172), .A(w62), .Cin(w164), .Cout(w178), .S(w182));   //: @(135, 860) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w52 = A[6]; //: TAP g72 @(-739,65) /sn:0 /R:1 /w:[ 1 46 45 ] /ss:1
  AND2 g153 (.in1(w92), .in2(w120), .out(w122));   //: @(-2605, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  FA g203 (.A(w36), .B(w141), .Cin(w135), .Cout(w149), .S(w150));   //: @(350, 680) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  AND2 g99 (.in1(w58), .in2(w64), .out(w70));   //: @(-1407, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  AND2 g98 (.in1(w58), .in2(w50), .out(w61));   //: @(-1354, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  //: joint g161 (w92) @(-2575, 325) /w:[ 2 -1 28 1 ]
  //: joint g182 (w109) @(-2892, 325) /w:[ 8 -1 7 22 ]
  FA g196 (.A(w25), .B(w11), .Cin(w143), .Cout(w147), .S(w141));   //: @(352, 499) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w69 = A[6]; //: TAP g96 @(-1204,65) /sn:0 /R:1 /w:[ 1 62 61 ] /ss:1
  //: joint g16 (w1) @(317, 317) /w:[ 4 -1 3 26 ]
  assign w128 = A[3]; //: TAP g189 @(-2913,65) /sn:0 /R:1 /w:[ 1 120 119 ] /ss:1
  //: joint g183 (w109) @(-2947, 325) /w:[ 6 -1 5 24 ]
  AND2 g152 (.in1(w92), .in2(w117), .out(w119));   //: @(-2554, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  AND2 g103 (.in1(w58), .in2(w83), .out(w85));   //: @(-1624, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  AND2 g122 (.in1(w75), .in2(w67), .out(w78));   //: @(-1822, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  FA g246 (.B(w240), .A(w133), .Cin(w245), .Cout(w251), .S(w252));   //: @(-207, 1502) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  assign w1 = B[0]; //: TAP g10 @(589,96) /sn:0 /R:1 /w:[ 15 2 1 ] /ss:1
  AND2 g78 (.in1(w41), .in2(w63), .out(w65));   //: @(-1104, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  //: joint g87 (w41) @(-1073, 323) /w:[ 6 -1 5 24 ]
  FA g212 (.B(w168), .A(w59), .Cin(w153), .Cout(w164), .S(w173));   //: @(202, 860) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g199 (.A(w34), .B(w20), .Cin(w155), .Cout(w159), .S(w160));   //: @(136, 499) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  AND2 g171 (.in1(w109), .in2(w115), .out(w121));   //: @(-2814, 359) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  AND2 g129 (.in1(w75), .in2(w103), .out(w105));   //: @(-2145, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  AND2 g27 (.in1(w7), .in2(w13), .out(w19));   //: @(-12, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  AND2 g32 (.in1(w7), .in2(w35), .out(w37));   //: @(-280, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  assign w115 = A[1]; //: TAP g187 @(-2805,65) /sn:0 /R:1 /w:[ 1 116 115 ] /ss:1
  AND2 g102 (.in1(w58), .in2(w80), .out(w82));   //: @(-1570, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  assign w100 = A[5]; //: TAP g143 @(-2080,65) /sn:0 /R:1 /w:[ 1 92 91 ] /ss:1
  assign w43 = A[3]; //: TAP g69 @(-574,65) /sn:0 /R:1 /w:[ 1 40 39 ] /ss:1
  FA g240 (.B(w232), .A(w122), .Cin(w239), .Cout(w243), .S(w244));   //: @(-282, 1322) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g244 (.B(w230), .A(w127), .Cin(w225), .Cout(w237), .S(w238));   //: @(-75, 1502) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  AND2 g9 (.in1(w1), .in2(w21), .out(w23));   //: @(179, 355) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  AND2 g57 (.in1(w56), .in2(w24), .out(w181));   //: @(-804, 355) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<0 ]
  assign w83 = A[5]; //: TAP g119 @(-1615,65) /sn:0 /R:1 /w:[ 1 76 75 ] /ss:1
  FA g245 (.B(w236), .A(w130), .Cin(w237), .Cout(w245), .S(w246));   //: @(-141, 1502) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  assign w97 = A[4]; //: TAP g142 @(-2026,65) /sn:0 /R:1 /w:[ 1 90 89 ] /ss:1
  //: joint g15 (w1) @(372, 317) /w:[ 6 -1 5 24 ]
  assign w49 = A[5]; //: TAP g71 @(-684,65) /sn:0 /R:1 /w:[ 1 44 43 ] /ss:1
  assign w84 = A[0]; //: TAP g162 @(-2284,65) /sn:0 /R:1 /w:[ 1 98 97 ] /ss:1
  //: joint g131 (w75) @(-1792, 323) /w:[ -1 14 13 16 ]
  assign w30 = A[1]; //: TAP g67 @(-464,65) /sn:0 /R:1 /w:[ 1 36 35 ] /ss:1
  assign w75 = B[5]; //: TAP g127 @(-1793,96) /sn:0 /R:1 /w:[ 15 12 11 ] /ss:1
  assign w13 = A[1]; //: TAP g43 @(-3,65) /sn:0 /R:1 /w:[ 1 20 19 ] /ss:1
  assign w106 = A[7]; //: TAP g145 @(-2188,65) /sn:0 /R:1 /w:[ 1 96 95 ] /ss:1
  //: joint g62 (w56) @(-550, 320) /w:[ 8 -1 7 22 ]
  assign w24 = A[7]; //: TAP g73 @(-793,65) /sn:0 /R:1 /w:[ 0 48 47 ] /ss:1
  //: joint g88 (w41) @(-1129, 323) /w:[ 4 -1 3 26 ]
  AND2 g104 (.in1(w58), .in2(w86), .out(w88));   //: @(-1678, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  assign w124 = A[2]; //: TAP g188 @(-2859,65) /sn:0 /R:1 /w:[ 1 118 117 ] /ss:1
  //: joint g180 (w109) @(-2785, 325) /w:[ 12 -1 11 18 ]
  assign w67 = A[0]; //: TAP g138 @(-1813,65) /sn:0 /R:1 /w:[ 1 82 81 ] /ss:1
  //: joint g42 (w7) @(-251, 324) /w:[ 2 -1 28 1 ]
  //: joint g63 (w56) @(-606, 320) /w:[ 6 -1 5 24 ]
  AND2 g175 (.in1(w109), .in2(w134), .out(w136));   //: @(-3030, 360) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  AND2 g74 (.in1(w41), .in2(w33), .out(w44));   //: @(-885, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  //: joint g109 (w58) @(-1430, 323) /w:[ 10 -1 9 20 ]
  HA g234 (.B(w194), .A(w95), .Cout(w162), .S(w185));   //: @(133, 1322) /sz:(40, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  //: joint g181 (w109) @(-2839, 325) /w:[ 10 -1 9 20 ]
  assign w120 = A[6]; //: TAP g168 @(-2594,65) /sn:0 /R:1 /w:[ 1 110 109 ] /ss:1
  //: joint g133 (w75) @(-1898, 323) /w:[ 10 -1 9 20 ]
  AND2 g5 (.in1(w1), .in2(w9), .out(w11));   //: @(398, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  AND2 g56 (.in1(w56), .in2(w52), .out(w54));   //: @(-749, 355) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  HA g194 (.A(w10), .B(w5), .Cout(w129), .S(w132));   //: @(496, 500) /sz:(40, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  AND2 g79 (.in1(w41), .in2(w66), .out(w68));   //: @(-1159, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  assign w66 = A[5]; //: TAP g95 @(-1150,65) /sn:0 /R:1 /w:[ 1 60 59 ] /ss:1
  assign w77 = A[3]; //: TAP g117 @(-1505,65) /sn:0 /R:1 /w:[ 1 72 71 ] /ss:1
  FA g215 (.B(w180), .A(w68), .Cin(w187), .Cout(w191), .S(w192));   //: @(0, 859) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w18 = A[6]; //: TAP g24 @(247,65) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  assign w4 = A[0]; //: TAP g36 @(50,65) /sn:0 /R:1 /w:[ 1 18 17 ] /ss:1
  //: joint g85 (w41) @(-966, 323) /w:[ 10 -1 9 20 ]
  assign w55 = A[2]; //: TAP g92 @(-986,65) /sn:0 /R:1 /w:[ 1 54 53 ] /ss:1
  FA g216 (.B(w184), .A(w71), .Cin(w191), .Cout(w195), .S(w196));   //: @(-67, 859) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w109 = B[7]; //: TAP g178 @(-2728,96) /sn:0 /R:1 /w:[ 15 16 15 ] /ss:1
  assign w103 = A[6]; //: TAP g144 @(-2136,65) /sn:0 /R:1 /w:[ 1 94 93 ] /ss:1
  AND2 g125 (.in1(w75), .in2(w94), .out(w96));   //: @(-1982, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  //: joint g60 (w56) @(-444, 320) /w:[ 12 -1 11 18 ]
  AND2 g81 (.in1(w41), .in2(w72), .out(w74));   //: @(-1268, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  AND2 g101 (.in1(w58), .in2(w77), .out(w79));   //: @(-1516, 357) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  HA g210 (.B(w150), .A(w44), .Cout(w57), .S(w118));   //: @(347, 861) /sz:(40, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  FA g214 (.B(w176), .A(w65), .Cin(w178), .Cout(w187), .S(w188));   //: @(66, 860) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g204 (.A(w42), .B(w152), .Cin(w149), .Cout(w157), .S(w158));   //: @(284, 680) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g185 (w109) @(-3053, 325) /w:[ 2 -1 28 1 ]
  AND2 g170 (.in1(w109), .in2(w101), .out(w112));   //: @(-2758, 359) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  assign w12 = A[4]; //: TAP g22 @(352,65) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  //: joint g35 (w7) @(71, 324) /w:[ -1 14 13 16 ]
  assign w26 = A[3]; //: TAP g45 @(-112,65) /sn:0 /R:1 /w:[ 1 24 23 ] /ss:1
  assign w46 = A[4]; //: TAP g70 @(-626,65) /sn:0 /R:1 /w:[ 1 42 41 ] /ss:1
  AND2 g126 (.in1(w75), .in2(w97), .out(w99));   //: @(-2035, 358) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  //: OUT g251 (S) @(132,1867) /sn:0 /w:[ 0 ]
  FA g209 (.A(w181), .B(w166), .Cin(w179), .Cout(w183), .S(w184));   //: @(-50, 677) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g184 (w109) @(-3001, 325) /w:[ 4 -1 3 26 ]
  assign w16 = A[0]; //: TAP g66 @(-413,65) /sn:0 /R:1 /w:[ 1 34 33 ] /ss:1
  assign w72 = A[7]; //: TAP g97 @(-1260,65) /sn:0 /R:1 /w:[ 1 64 63 ] /ss:1
  assign w50 = A[0]; //: TAP g114 @(-1343,65) /sn:0 /R:1 /w:[ 1 66 65 ] /ss:1
  assign w86 = A[6]; //: TAP g120 @(-1667,65) /sn:0 /R:1 /w:[ 1 78 77 ] /ss:1
  FA g235 (.B(w206), .A(w104), .Cin(w162), .Cout(w209), .S(w210));   //: @(66, 1321) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g12 (w1) @(535, 317) /w:[ 12 -1 11 18 ]
  assign w0 = A[0]; //: TAP g18 @(569,65) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  HA g226 (.B(w177), .A(w78), .Cout(w148), .S(w161));   //: @(205, 1160) /sz:(40, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  FA g229 (.B(w204), .A(w96), .Cin(w205), .Cout(w213), .S(w214));   //: @(-2, 1159) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w134 = A[5]; //: TAP g191 @(-3019,65) /sn:0 /R:1 /w:[ 1 124 123 ] /ss:1
  assign w107 = A[2]; //: TAP g164 @(-2388,65) /sn:0 /R:1 /w:[ 1 102 101 ] /ss:1
  AND2 g30 (.in1(w7), .in2(w29), .out(w31));   //: @(-173, 356) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  //: joint g108 (w58) @(-1377, 323) /w:[ 12 -1 11 18 ]
  FA g219 (.B(w173), .A(w70), .Cin(w145), .Cout(w174), .S(w177));   //: @(201, 1001) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g239 (.B(w228), .A(w119), .Cin(w235), .Cout(w239), .S(w240));   //: @(-214, 1323) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g134 (w75) @(-1951, 323) /w:[ 8 -1 7 22 ]
  assign w80 = A[4]; //: TAP g118 @(-1561,65) /sn:0 /R:1 /w:[ 1 74 73 ] /ss:1
  HA g242 (.B(w210), .A(w112), .Cout(w186), .S(w201));   //: @(64, 1501) /sz:(40, 54) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FS
module FS(D, Bout, Bin, B, A);
//: interface  /sz:(53, 64) /bd:[ Ti0>A(13/53) Ti1>B(39/53) Ri0>Bin(28/64) Lo0<Bout(27/64) Bo0<D(25/53) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(242,272)(138,272)(138,111){1}
//: {2}(140,109)(158,109){3}
//: {4}(136,109)(123,109){5}
input A;    //: /sn:0 {0}(164,242)(146,242)(146,93){1}
//: {2}(148,91)(158,91){3}
//: {4}(144,91)(123,91){5}
output Bout;    //: /sn:0 {0}(593,248)(530,248)(530,248)(547,248){1}
output D;    //: /sn:0 {0}(402,125)(326,125){1}
input Bin;    //: /sn:0 {0}(350,208)(235,208)(235,140){1}
//: {2}(237,138)(256,138)(256,126)(269,126){3}
//: {4}(233,138)(197,138){5}
wire w6;    //: /sn:0 {0}(505,249)(473,249){1}
wire w7;    //: /sn:0 {0}(431,239)(407,239)(407,197)(392,197){1}
wire w4;    //: /sn:0 {0}(431,261)(299,261)(299,261)(284,261){1}
wire w3;    //: /sn:0 {0}(350,188)(334,188)(334,177)(319,177){1}
wire w1;    //: /sn:0 {0}(242,252)(221,252)(221,241)(206,241){1}
wire w2;    //: /sn:0 {0}(277,178)(250,178)(250,110){1}
//: {2}(252,108)(269,108){3}
//: {4}(248,108)(215,108){5}
//: enddecls

  //: OUT g4 (D) @(399,125) /sn:0 /w:[ 0 ]
  //: joint g8 (A) @(146, 91) /w:[ 2 -1 4 1 ]
  //: OUT g3 (Bout) @(590,248) /sn:0 /w:[ 0 ]
  //: joint g13 (w2) @(250, 108) /w:[ 2 -1 4 1 ]
  //: IN g2 (Bin) @(195,138) /sn:0 /w:[ 5 ]
  //: IN g1 (B) @(121,109) /sn:0 /w:[ 5 ]
  INV1 g11 (.in(w2), .out(w3));   //: @(278, 157) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  INV1 g16 (.in(w6), .out(Bout));   //: @(506, 228) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  //: joint g10 (B) @(138, 109) /w:[ 2 -1 4 1 ]
  EXOR2 g6 (.b(Bin), .a(w2), .out(D));   //: @(270, 98) /sz:(55, 42) /sn:0 /p:[ Li0>3 Li1>3 Ro0<1 ]
  INV1 g7 (.in(A), .out(w1));   //: @(165, 221) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  AND2 g9 (.in2(B), .in1(w1), .out(w4));   //: @(243, 242) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  NOR2 g15 (.in2(w4), .in1(w7), .out(w6));   //: @(432, 231) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  EXOR2 g5 (.b(B), .a(A), .out(w2));   //: @(159, 81) /sz:(55, 42) /sn:0 /p:[ Li0>3 Li1>3 Ro0<5 ]
  //: joint g14 (Bin) @(235, 138) /w:[ 2 -1 4 1 ]
  //: IN g0 (A) @(121,91) /sn:0 /w:[ 5 ]
  AND2 g12 (.in2(Bin), .in1(w3), .out(w7));   //: @(351, 178) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX2
module MUX2(out, c, in0, in1);
//: interface  /sz:(40, 42) /bd:[ Li0>in0(9/42) Li1>in1(28/42) Bi0>c(23/40) Ro0<out(18/42) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output out;    //: /sn:0 {0}(472,139)(396,139)(396,155)(381,155){1}
input in0;    //: /sn:0 {0}(78,83)(210,83)(210,88)(225,88){1}
input in1;    //: /sn:0 {0}(75,208)(206,208)(206,207)(221,207){1}
input c;    //: /sn:0 {0}(158,302)(158,229){1}
//: {2}(160,227)(221,227){3}
//: {4}(158,225)(158,196)(153,196)(153,183){5}
wire w1;    //: /sn:0 {0}(152,141)(152,108)(225,108){1}
wire w2;    //: /sn:0 {0}(267,96)(324,96)(324,147)(339,147){1}
wire w5;    //: /sn:0 {0}(263,215)(324,215)(324,167)(339,167){1}
//: enddecls

  //: OUT g8 (out) @(469,139) /sn:0 /w:[ 0 ]
  //: IN g4 (c) @(158,304) /sn:0 /R:1 /w:[ 0 ]
  INV1 g3 (.in(c), .out(w1));   //: @(132, 142) /sz:(40, 40) /R:1 /sn:0 /p:[ Bi0>5 To0<0 ]
  NAND2 g2 (.in2(w5), .in1(w2), .out(out));   //: @(340, 137) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 ]
  NAND2 g1 (.in2(c), .in1(in1), .out(w5));   //: @(222, 197) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]
  //: IN g6 (in0) @(76,83) /sn:0 /w:[ 0 ]
  //: IN g7 (in1) @(73,208) /sn:0 /w:[ 0 ]
  //: joint g5 (c) @(158, 227) /w:[ 2 4 -1 1 ]
  NAND2 g0 (.in2(w1), .in1(in0), .out(w2));   //: @(226, 78) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin INV1
module INV1(in, out);
//: interface  /sz:(40, 40) /bd:[ Li0>in(21/40) Ro0<out(20/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w6;    //: /sn:0 {0}(320,88)(320,142)(320,142)(320,123){1}
input in;    //: /sn:0 {0}(235,162)(289,162){1}
//: {2}(291,160)(291,131)(306,131){3}
//: {4}(291,164)(291,200)(306,200){5}
output out;    //: /sn:0 {0}(320,192)(320,164){1}
//: {2}(322,162)(332,162)(332,162)(373,162){3}
//: {4}(320,160)(320,140){5}
supply0 w3;    //: /sn:0 {0}(320,209)(320,215)(320,215)(320,230){1}
//: enddecls

  //: IN g4 (in) @(233,162) /sn:0 /w:[ 0 ]
  //: VDD g3 (w6) @(331,88) /sn:0 /w:[ 0 ]
  //: GROUND g2 (w3) @(320,236) /sn:0 /w:[ 1 ]
  _GGNMOS #(2, 1) g1 (.Z(out), .S(w3), .G(in));   //: @(314,200) /sn:0 /w:[ 0 0 5 ]
  //: joint g6 (in) @(291, 162) /w:[ -1 2 1 4 ]
  //: joint g7 (out) @(320, 162) /w:[ 2 4 -1 1 ]
  //: OUT g5 (out) @(370,162) /sn:0 /w:[ 3 ]
  _GGPMOS #(2, 1) g0 (.Z(out), .S(w6), .G(in));   //: @(314,131) /sn:0 /w:[ 5 1 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin Div8b
module Div8b(D, B, A, R);
//: interface  /sz:(80, 64) /bd:[ Li0>B[7:0](46/64) Li1>A[7:0](16/64) Bo0<R[7:0](60/80) Bo1<D[7:0](20/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply0 w32;    //: /sn:0 {0}(798,214)(798,232)(743,232){1}
input [7:0] A;    //: /sn:0 {0}(#:58,82)(699,82){1}
//: {2}(700,82)(928,82){3}
//: {4}(929,82)(1362,82)(1362,359){5}
//: {6}(1362,360)(1362,583){7}
//: {8}(1362,584)(1362,739){9}
//: {10}(1362,740)(1362,1226){11}
//: {12}(1362,1227)(1362,2384){13}
//: {14}(1362,2385)(1362,2819){15}
//: {16}(1362,2820)(1362,2834){17}
supply0 w225;    //: /sn:0 {0}(1304,2661)(1304,2682)(1282,2682){1}
supply0 w126;    //: /sn:0 {0}(1009,1427)(1009,1447)(994,1447){1}
supply0 w37;    //: /sn:0 {0}(894,1021)(894,1036)(877,1036){1}
supply0 w128;    //: /sn:0 {0}(1084,1865)(1084,1879)(1063,1879){1}
supply0 w258;    //: /sn:0 {0}(1410,3090)(1410,3106)(1394,3106){1}
supply0 w192;    //: /sn:0 {0}(1186,2253)(1186,2275)(1170,2275){1}
output [7:0] D;    //: /sn:0 {0}(238,3436)(194,3436)(#:194,3418){1}
input [7:0] B;    //: /sn:0 {0}(#:58,129)(168,129){1}
//: {2}(169,129)(253,129){3}
//: {4}(254,129)(334,129){5}
//: {6}(335,129)(418,129){7}
//: {8}(419,129)(495,129){9}
//: {10}(496,129)(576,129){11}
//: {12}(577,129)(651,129){13}
//: {14}(652,129)(727,129){15}
//: {16}(728,129)(826,129)(826,542){17}
//: {18}(824,544)(807,544){19}
//: {20}(806,544)(738,544){21}
//: {22}(737,544)(658,544){23}
//: {24}(657,544)(573,544){25}
//: {26}(572,544)(487,544){27}
//: {28}(486,544)(407,544){29}
//: {30}(406,544)(326,544){31}
//: {32}(325,544)(242,544){33}
//: {34}(241,544)(115,544)(115,967){35}
//: {36}(117,969)(259,969){37}
//: {38}(260,969)(346,969){39}
//: {40}(347,969)(430,969){41}
//: {42}(431,969)(511,969){43}
//: {44}(512,969)(592,969){45}
//: {46}(593,969)(680,969){47}
//: {48}(681,969)(772,969){49}
//: {50}(773,969)(860,969){51}
//: {52}(861,969)(1039,969)(1039,1372){53}
//: {54}(1037,1374)(978,1374){55}
//: {56}(977,1374)(890,1374){57}
//: {58}(889,1374)(796,1374){59}
//: {60}(795,1374)(706,1374){61}
//: {62}(705,1374)(618,1374){63}
//: {64}(617,1374)(530,1374){65}
//: {66}(529,1374)(447,1374){67}
//: {68}(446,1374)(367,1374){69}
//: {70}(366,1374)(279,1374)(279,1804){71}
//: {72}(281,1806)(473,1806){73}
//: {74}(474,1806)(553,1806){75}
//: {76}(554,1806)(638,1806){77}
//: {78}(639,1806)(719,1806){79}
//: {80}(720,1806)(783,1806){81}
//: {82}(784,1806)(881,1806){83}
//: {84}(882,1806)(967,1806){85}
//: {86}(968,1806)(1048,1806){87}
//: {88}(1049,1806)(1086,1806){89}
//: {90}(279,1808)(279,2206)(281,2206){91}
//: {92}(285,2206)(576,2206){93}
//: {94}(577,2206)(658,2206){95}
//: {96}(659,2206)(742,2206){97}
//: {98}(743,2206)(820,2206){99}
//: {100}(821,2206)(903,2206){101}
//: {102}(904,2206)(988,2206){103}
//: {104}(989,2206)(1068,2206){105}
//: {106}(1069,2206)(1153,2206){107}
//: {108}(1154,2206)(1194,2206){109}
//: {110}(283,2208)(283,2607)(300,2607){111}
//: {112}(304,2607)(680,2607){113}
//: {114}(681,2607)(763,2607){115}
//: {116}(764,2607)(843,2607){117}
//: {118}(844,2607)(925,2607){119}
//: {120}(926,2607)(1010,2607){121}
//: {122}(1011,2607)(1090,2607){123}
//: {124}(1091,2607)(1175,2607){125}
//: {126}(1176,2607)(1265,2607){127}
//: {128}(1266,2607)(1297,2607){129}
//: {130}(302,2609)(302,3027)(785,3027){131}
//: {132}(786,3027)(865,3027){133}
//: {134}(866,3027)(948,3027){135}
//: {136}(949,3027)(1032,3027){137}
//: {138}(1033,3027)(1112,3027){139}
//: {140}(1113,3027)(1198,3027){141}
//: {142}(1199,3027)(1287,3027){143}
//: {144}(1288,3027)(1378,3027){145}
//: {146}(1379,3027)(1414,3027){147}
//: {148}(1039,1376)(1039,1387){149}
//: {150}(115,971)(115,978){151}
//: {152}(826,546)(826,550){153}
output [7:0] R;    //: /sn:0 {0}(1112,3623)(1076,3623)(#:1076,3581){1}
supply0 w31;    //: /sn:0 {0}(658,432)(658,314)(600,314)(600,182)(625,182){1}
//: {2}(627,180)(627,174)(552,174){3}
//: {4}(550,172)(550,146)(529,146)(529,310)(578,310)(578,409){5}
//: {6}(548,174)(475,174){7}
//: {8}(471,174)(397,174){9}
//: {10}(393,174)(315,174){11}
//: {12}(313,172)(313,157)(288,157)(288,305)(324,305)(324,338){13}
//: {14}(311,174)(232,174){15}
//: {16}(230,172)(230,162)(201,162)(201,297)(242,297)(242,315){17}
//: {18}(228,174)(145,174){19}
//: {20}(141,174)(113,174){21}
//: {22}(143,176)(143,196){23}
//: {24}(230,176)(230,197){25}
//: {26}(313,176)(313,198){27}
//: {28}(395,176)(395,184)(393,184)(393,187){29}
//: {30}(391,189)(365,189)(365,304)(412,304)(412,360){31}
//: {32}(393,191)(393,199){33}
//: {34}(473,176)(473,184)(472,184)(472,187){35}
//: {36}(470,189)(444,189)(444,305)(496,305)(496,384){37}
//: {38}(472,191)(472,200){39}
//: {40}(550,176)(550,201){41}
//: {42}(627,184)(627,202){43}
supply0 w59;    //: /sn:0 {0}(880,595)(880,608)(850,608){1}
wire w270;    //: /sn:0 {0}(1041,3575)(1041,3556)(783,3556)(783,3251){1}
wire w96;    //: /sn:0 {0}(507,1199)(507,1119)(460,1119)(460,989)(487,989){1}
//: {2}(489,987)(489,956)(575,956)(575,864){3}
//: {4}(489,991)(489,1004){5}
wire w73;    //: /sn:0 {0}(431,973)(431,1003){1}
wire w45;    //: /sn:0 {0}(416,768)(416,721)(393,721)(393,640){1}
wire w160;    //: /sn:0 {0}(729,2413)(729,2350)(688,2350)(688,2228)(715,2228){1}
//: {2}(717,2226)(717,2079){3}
//: {4}(717,2230)(717,2241){5}
wire w244;    //: /sn:0 {0}(935,3138)(935,3170)(954,3170)(954,3261){1}
wire w56;    //: /sn:0 {0}(812,903)(812,675)(774,675)(774,560)(817,560)(817,562){1}
//: {2}(819,564)(929,564)(929,86){3}
//: {4}(815,564)(809,564)(809,579){5}
wire w16;    //: /sn:0 {0}(496,133)(496,141)(498,141)(498,200){1}
wire w218;    //: /sn:0 {0}(1137,2680)(1119,2680)(1119,2680)(1107,2680){1}
wire w266;    //: /sn:0 {0}(169,3412)(169,3383)(63,3383)(63,3307){1}
wire w89;    //: /sn:0 {0}(822,1035)(801,1035)(801,1036)(789,1036){1}
wire w81;    //: /sn:0 {0}(681,973)(681,981)(682,981)(682,1006){1}
wire w19;    //: /sn:0 {0}(536,229)(513,229){1}
wire w4;    //: /sn:0 {0}(155,277)(155,262){1}
wire w183;    //: /sn:0 {0}(990,2244)(990,2218)(989,2218)(989,2210){1}
wire w0;    //: /sn:0 {0}(169,133)(169,196){1}
wire w151;    //: /sn:0 {0}(706,1912)(706,1942)(726,1942)(726,2037){1}
wire w120;    //: /sn:0 {0}(978,1378)(978,1386)(979,1386)(979,1418){1}
wire w233;    //: /sn:0 {0}(1100,3319)(1100,3196)(1060,3196)(1060,3059)(1086,3059){1}
//: {2}(1088,3057)(1088,2945){3}
//: {4}(1088,3061)(1088,3074){5}
wire w240;    //: /sn:0 {0}(949,3072)(949,3031){1}
wire w111;    //: /sn:0 {0}(706,1378)(706,1386)(708,1386)(708,1415){1}
wire w104;    //: /sn:0 {0}(162,3265)(162,3251)(157,3251)(157,1585){1}
//: {2}(159,1583)(361,1583){3}
//: {4}(365,1583)(420,1583){5}
//: {6}(363,1585)(363,1610){7}
//: {8}(365,1612)(507,1612){9}
//: {10}(363,1614)(363,1646){11}
//: {12}(365,1648)(595,1648){13}
//: {14}(363,1650)(363,1675){15}
//: {16}(365,1677)(574,1677)(574,1677)(684,1677){17}
//: {18}(363,1679)(363,1704){19}
//: {20}(365,1706)(773,1706){21}
//: {22}(363,1708)(363,1734){23}
//: {24}(365,1736)(868,1736){25}
//: {26}(363,1738)(363,1764)(947,1764){27}
//: {28}(157,1581)(157,1439)(329,1439){29}
wire w168;    //: /sn:0 {0}(976,2499)(976,2378)(935,2378)(935,2226)(962,2226){1}
//: {2}(964,2224)(964,2153){3}
//: {4}(964,2228)(964,2244){5}
wire w171;    //: /sn:0 {0}(562,2305)(562,2320){1}
wire w237;    //: /sn:0 {0}(773,3136)(773,3165)(792,3165)(792,3209){1}
wire w119;    //: /sn:0 {0}(851,1445)(814,1445){1}
wire w67;    //: /sn:0 {0}(589,1224)(589,1113)(541,1113)(541,994)(567,994){1}
//: {2}(569,992)(569,932)(661,932)(661,892){3}
//: {4}(569,996)(569,1005){5}
wire w54;    //: /sn:0 {0}(644,643)(644,671)(670,671)(670,850){1}
wire w90;    //: /sn:0 {0}(850,1295)(850,1120)(808,1120)(808,992)(834,992){1}
//: {2}(836,990)(836,981)(992,981)(992,360)(1357,360){3}
//: {4}(836,994)(836,1007){5}
wire w176;    //: /sn:0 {0}(783,2270)(770,2270)(770,2270)(758,2270){1}
wire w167;    //: /sn:0 {0}(1034,1916)(1034,1943)(1053,1943)(1053,2135){1}
wire w124;    //: /sn:0 {0}(877,1483)(877,1512)(902,1512)(902,1712){1}
wire w23;    //: /sn:0 {0}(613,230)(599,230)(599,230)(591,230){1}
wire w20;    //: /sn:0 {0}(577,133)(577,141)(576,141)(576,201){1}
wire w174;    //: /sn:0 {0}(743,2241)(743,2210){1}
wire w272;    //: /sn:0 {0}(1061,3575)(1061,3539)(945,3539)(945,3303){1}
wire w108;    //: /sn:0 {0}(618,1378)(618,1386)(619,1386)(619,1414){1}
wire w223;    //: /sn:0 {0}(1163,2718)(1163,2749)(1182,2749)(1182,2930){1}
wire w125;    //: /sn:0 {0}(474,1810)(474,1818)(473,1818)(473,1843){1}
wire w103;    //: /sn:0 {0}(883,1712)(883,1590)(831,1590)(831,1401)(863,1401){1}
//: {2}(865,1399)(865,1348)(860,1348)(860,1337){3}
//: {4}(865,1403)(865,1417){5}
wire w8;    //: /sn:0 {0}(335,133)(335,141)(339,141)(339,198){1}
wire w71;    //: /sn:0 {0}(112,3265)(112,1167){1}
//: {2}(114,1165)(140,1165){3}
//: {4}(144,1165)(318,1165){5}
//: {6}(142,1167)(142,1190){7}
//: {8}(144,1192)(403,1192){9}
//: {10}(142,1194)(142,1221){11}
//: {12}(144,1223)(492,1223){13}
//: {14}(142,1225)(142,1246){15}
//: {16}(144,1248)(574,1248){17}
//: {18}(142,1250)(142,1269){19}
//: {20}(144,1271)(660,1271){21}
//: {22}(142,1273)(142,1292){23}
//: {24}(144,1294)(752,1294){25}
//: {26}(142,1296)(142,1319)(835,1319){27}
//: {28}(112,1163)(112,1029)(222,1029){29}
wire w202;    //: /sn:0 {0}(913,2845)(913,2777)(871,2777)(871,2636)(899,2636){1}
//: {2}(901,2634)(901,2516){3}
//: {4}(901,2638)(901,2649){5}
wire w238;    //: /sn:0 {0}(867,3071)(867,3039)(866,3039)(866,3031){1}
wire w17;    //: /sn:0 {0}(405,265)(405,293)(431,293)(431,360){1}
wire w84;    //: /sn:0 {0}(773,973)(773,981)(774,981)(774,1007){1}
wire w53;    //: /sn:0 {0}(807,548)(807,556)(835,556)(835,579){1}
wire w263;    //: /sn:0 {0}(199,3412)(199,3323)(218,3323)(218,3308){1}
wire w255;    //: /sn:0 {0}(1379,3077)(1379,3031){1}
wire w211;    //: /sn:0 {0}(831,2714)(831,2746)(850,2746)(850,2816){1}
wire w113;    //: /sn:0 {0}(668,1443)(634,1443){1}
wire w44;    //: /sn:0 {0}(573,548)(573,556)(574,556)(574,576){1}
wire w2;    //: /sn:0 {0}(216,225)(173,225)(173,225)(184,225){1}
wire w115;    //: /sn:0 {0}(605,1480)(605,1508)(629,1508)(629,1624){1}
wire w83;    //: /sn:0 {0}(642,1034)(610,1034){1}
wire w77;    //: /sn:0 {0}(475,1032)(459,1032)(459,1032)(446,1032){1}
wire w274;    //: /sn:0 {0}(1081,3575)(1081,3527)(1110,3527)(1110,3361){1}
wire w262;    //: /sn:0 {0}(209,3412)(209,3376)(275,3376)(275,3308){1}
wire w224;    //: /sn:0 {0}(1365,3387)(1365,3204)(1320,3204)(1320,3058)(1351,3058){1}
//: {2}(1353,3056)(1353,2820)(1357,2820){3}
//: {4}(1353,3060)(1353,3077){5}
wire w10;    //: /sn:0 {0}(286,601)(264,601)(264,601)(256,601){1}
wire w275;    //: /sn:0 {0}(1091,3575)(1091,3541)(1195,3541)(1195,3383){1}
wire w273;    //: /sn:0 {0}(1071,3575)(1071,3526)(1030,3526)(1030,3332){1}
wire w190;    //: /sn:0 {0}(1056,2311)(1056,2339)(1075,2339)(1075,2527){1}
wire w95;    //: /sn:0 {0}(343,1183)(343,1396)(343,1396)(343,1411){1}
wire w52;    //: /sn:0 {0}(701,606)(681,606)(681,606)(673,606){1}
wire w188;    //: /sn:0 {0}(1115,2274)(1100,2274)(1100,2274)(1085,2274){1}
wire w142;    //: /sn:0 {0}(639,1810)(639,1818)(638,1818)(638,1845){1}
wire w155;    //: /sn:0 {0}(787,1913)(787,1956)(806,1956)(806,2062){1}
wire w178;    //: /sn:0 {0}(729,2307)(729,2336)(748,2336)(748,2413){1}
wire w187;    //: /sn:0 {0}(976,2310)(976,2339)(995,2339)(995,2499){1}
wire w50;    //: /sn:0 {0}(738,548)(738,556)(741,556)(741,578){1}
wire w6;    //: /sn:0 {0}(326,548)(326,573){1}
wire w7;    //: /sn:0 {0}(299,226)(282,226)(282,226)(271,226){1}
wire w99;    //: /sn:0 {0}(522,1588)(522,1524)(474,1524)(474,1397)(502,1397){1}
//: {2}(504,1395)(504,1252)(517,1252)(517,1241){3}
//: {4}(504,1399)(504,1413){5}
wire w61;    //: /sn:0 {0}(347,973)(347,1002){1}
wire w135;    //: /sn:0 {0}(869,2088)(869,2005)(826,2005)(826,1831)(855,1831){1}
//: {2}(857,1829)(857,1765)(893,1765)(893,1754){3}
//: {4}(857,1833)(857,1848){5}
wire w153;    //: /sn:0 {0}(843,1876)(824,1876)(824,1876)(816,1876){1}
wire w216;    //: /sn:0 {0}(1092,2651)(1092,2619)(1091,2619)(1091,2611){1}
wire w106;    //: /sn:0 {0}(530,1378)(530,1413){1}
wire w69;    //: /sn:0 {0}(675,1247)(675,1124)(623,1124)(623,994)(654,994){1}
//: {2}(656,992)(656,941)(748,941)(748,918){3}
//: {4}(656,996)(656,1006){5}
wire w51;    //: /sn:0 {0}(584,822)(584,661)(560,661)(560,642){1}
wire w207;    //: /sn:0 {0}(845,2648)(845,2619)(844,2619)(844,2611){1}
wire w213;    //: /sn:0 {0}(1012,2650)(1012,2619)(1011,2619)(1011,2611){1}
wire w239;    //: /sn:0 {0}(909,3100)(892,3100)(892,3100)(882,3100){1}
wire w271;    //: /sn:0 {0}(1051,3575)(1051,3547)(863,3547)(863,3276){1}
wire w66;    //: /sn:0 {0}(418,1168)(418,1103)(374,1103)(374,990)(403,990){1}
//: {2}(405,988)(405,942)(490,942)(490,838){3}
//: {4}(405,992)(405,1003){5}
wire w177;    //: /sn:0 {0}(823,2242)(823,2218)(821,2218)(821,2210){1}
wire w34;    //: /sn:0 {0}(565,822)(565,708)(517,708)(517,563)(546,563){1}
//: {2}(548,561)(548,505)(588,505)(588,451){3}
//: {4}(548,565)(548,576){5}
wire w234;    //: /sn:0 {0}(1185,3341)(1185,3189)(1144,3189)(1144,3061)(1171,3061){1}
//: {2}(1173,3059)(1173,2972){3}
//: {4}(1173,3063)(1173,3075){5}
wire w102;    //: /sn:0 {0}(788,1682)(788,1558)(740,1558)(740,1402)(771,1402){1}
//: {2}(773,1400)(773,1323)(777,1323)(777,1312){3}
//: {4}(773,1404)(773,1416){5}
wire w87;    //: /sn:0 {0}(861,973)(861,981)(862,981)(862,1007){1}
wire w43;    //: /sn:0 {0}(448,603)(431,603)(431,603)(422,603){1}
wire w157;    //: /sn:0 {0}(928,1877)(909,1877)(909,1877)(898,1877){1}
wire w254;    //: /sn:0 {0}(1339,3105)(1304,3105){1}
wire w58;    //: /sn:0 {0}(260,973)(260,981)(262,981)(262,1001){1}
wire w28;    //: /sn:0 {0}(728,133)(728,203){1}
wire w130;    //: /sn:0 {0}(445,1601)(445,1828)(447,1828)(447,1843){1}
wire w169;    //: /sn:0 {0}(1056,2527)(1056,2373)(1017,2373)(1017,2230)(1042,2230){1}
//: {2}(1044,2228)(1044,2177){3}
//: {4}(1044,2232)(1044,2245){5}
wire w132;    //: /sn:0 {0}(541,1910)(541,1926)(560,1926)(560,1984){1}
wire w184;    //: /sn:0 {0}(891,2309)(891,2341)(910,2341)(910,2474){1}
wire w25;    //: /sn:0 {0}(562,267)(562,291)(597,291)(597,409){1}
wire w65;    //: /sn:0 {0}(333,1141)(333,1101)(291,1101)(291,988)(319,988){1}
//: {2}(321,986)(321,939)(407,939)(407,810){3}
//: {4}(321,990)(321,1002){5}
wire w210;    //: /sn:0 {0}(927,2649)(927,2619)(926,2619)(926,2611){1}
wire w121;    //: /sn:0 {0}(785,1482)(785,1514)(807,1514)(807,1682){1}
wire w92;    //: /sn:0 {0}(409,1440)(386,1440)(386,1440)(384,1440){1}
wire w40;    //: /sn:0 {0}(367,602)(348,602)(348,602)(341,602){1}
wire w30;    //: /sn:0 {0}(734,457)(734,344)(684,344)(684,185)(700,185){1}
//: {2}(702,183)(702,90)(700,90)(700,86){3}
//: {4}(702,187)(702,203){5}
wire w162;    //: /sn:0 {0}(1049,1810)(1049,1818)(1048,1818)(1048,1850){1}
wire w217;    //: /sn:0 {0}(998,2716)(998,2742)(1017,2742)(1017,2875){1}
wire w149;    //: /sn:0 {0}(761,1875)(742,1875)(742,1875)(735,1875){1}
wire w146;    //: /sn:0 {0}(720,1810)(720,1846){1}
wire w222;    //: /sn:0 {0}(1267,2653)(1267,2619)(1266,2619)(1266,2611){1}
wire w165;    //: /sn:0 {0}(809,2445)(809,2371)(770,2371)(770,2231)(795,2231){1}
//: {2}(797,2229)(797,2104){3}
//: {4}(797,2233)(797,2242){5}
wire w248;    //: /sn:0 {0}(1129,3103)(1144,3103)(1144,3103)(1159,3103){1}
wire w139;    //: /sn:0 {0}(554,1810)(554,1818)(555,1818)(555,1844){1}
wire w136;    //: /sn:0 {0}(954,2111)(954,1985)(912,1985)(912,1834)(940,1834){1}
//: {2}(942,1832)(942,1793)(972,1793)(972,1782){3}
//: {4}(942,1836)(942,1849){5}
wire w49;    //: /sn:0 {0}(618,605)(598,605)(598,605)(589,605){1}
wire w57;    //: /sn:0 {0}(727,644)(727,674)(757,674)(757,876){1}
wire w173;    //: /sn:0 {0}(703,2269)(683,2269)(683,2269)(675,2269){1}
wire w105;    //: /sn:0 {0}(355,1492)(355,1477){1}
wire w148;    //: /sn:0 {0}(620,2268)(588,2268)(588,2268)(591,2268){1}
wire w252;    //: /sn:0 {0}(1289,3076)(1289,3039)(1288,3039)(1288,3031){1}
wire w186;    //: /sn:0 {0}(1070,2245)(1070,2218)(1069,2218)(1069,2210){1}
wire w72;    //: /sn:0 {0}(248,1082)(248,1067){1}
wire w94;    //: /sn:0 {0}(848,1073)(848,1097)(869,1097)(869,1295){1}
wire w33;    //: /sn:0 {0}(714,269)(714,292)(753,292)(753,457){1}
wire w191;    //: /sn:0 {0}(1253,2962)(1253,2825)(1211,2825)(1211,2641)(1239,2641){1}
//: {2}(1241,2639)(1241,2385)(1357,2385){3}
//: {4}(1241,2643)(1241,2653){5}
wire w107;    //: /sn:0 {0}(490,1441)(473,1441)(473,1441)(464,1441){1}
wire w145;    //: /sn:0 {0}(680,1874)(662,1874)(662,1874)(653,1874){1}
wire w9;    //: /sn:0 {0}(242,263)(242,280)(261,280)(261,315){1}
wire w79;    //: /sn:0 {0}(417,1069)(417,1096)(437,1096)(437,1168){1}
wire w219;    //: /sn:0 {0}(1177,2652)(1177,2619)(1176,2619)(1176,2611){1}
wire w39;    //: /sn:0 {0}(407,548)(407,574){1}
wire w55;    //: /sn:0 {0}(756,607)(795,607){1}
wire w201;    //: /sn:0 {0}(330,3266)(330,3029)(325,3029)(325,2792){1}
//: {2}(327,2790)(335,2790)(335,2791)(548,2791){3}
//: {4}(552,2791)(736,2791){5}
//: {6}(550,2793)(550,2838){7}
//: {8}(552,2840)(816,2840){9}
//: {10}(550,2842)(550,2867){11}
//: {12}(552,2869)(898,2869){13}
//: {14}(550,2871)(550,2897){15}
//: {16}(552,2899)(983,2899){17}
//: {18}(550,2901)(550,2925){19}
//: {20}(552,2927)(1063,2927){21}
//: {22}(550,2929)(550,2952){23}
//: {24}(552,2954)(1148,2954){25}
//: {26}(550,2956)(550,2986)(1238,2986){27}
//: {28}(325,2788)(325,2674)(642,2674){29}
wire w232;    //: /sn:0 {0}(1020,3290)(1020,3195)(979,3195)(979,3060)(1006,3060){1}
//: {2}(1008,3058)(1008,2917){3}
//: {4}(1008,3062)(1008,3073){5}
wire w122;    //: /sn:0 {0}(939,1446)(913,1446)(913,1446)(906,1446){1}
wire w134;    //: /sn:0 {0}(787,2062)(787,1965)(755,1965)(755,1820)(785,1820)(785,1828){1}
//: {2}(787,1830)(798,1830)(798,1724){3}
//: {4}(783,1830)(775,1830)(775,1847){5}
wire w166;    //: /sn:0 {0}(891,2474)(891,2345)(850,2345)(850,2226)(877,2226){1}
//: {2}(879,2224)(879,2130){3}
//: {4}(879,2228)(879,2243){5}
wire w203;    //: /sn:0 {0}(668,2712)(668,2727){1}
wire w214;    //: /sn:0 {0}(913,2715)(913,2749)(932,2749)(932,2845){1}
wire w14;    //: /sn:0 {0}(215,572)(215,462)(252,462)(252,357){1}
wire w141;    //: /sn:0 {0}(598,1873)(577,1873)(577,1873)(570,1873){1}
wire w220;    //: /sn:0 {0}(1078,2717)(1078,2743)(1097,2743)(1097,2903){1}
wire w179;    //: /sn:0 {0}(865,2271)(844,2271)(844,2271)(838,2271){1}
wire w38;    //: /sn:0 {0}(227,652)(227,638){1}
wire w195;    //: /sn:0 {0}(725,2675)(712,2675)(712,2675)(697,2675){1}
wire w250;    //: /sn:0 {0}(1100,3140)(1100,3168)(1119,3168)(1119,3319){1}
wire w152;    //: /sn:0 {0}(550,2239)(550,2042)(551,2042)(551,2026){1}
wire w180;    //: /sn:0 {0}(905,2243)(905,2218)(904,2218)(904,2210){1}
wire w182;    //: /sn:0 {0}(950,2272)(933,2272)(933,2272)(920,2272){1}
wire w3;    //: /sn:0 {0}(719,481)(206,481)(206,458){1}
//: {2}(208,456)(643,456){3}
//: {4}(206,454)(206,435){5}
//: {6}(208,433)(563,433){7}
//: {8}(206,431)(206,410){9}
//: {10}(208,408)(481,408){11}
//: {12}(206,406)(206,386){13}
//: {14}(208,384)(397,384){15}
//: {16}(206,382)(206,364){17}
//: {18}(208,362)(309,362){19}
//: {20}(206,360)(206,335){21}
//: {22}(208,333)(227,333){23}
//: {24}(204,333)(44,333){25}
//: {26}(42,331)(42,224)(129,224){27}
//: {28}(42,335)(42,3250)(8,3250)(8,3265){29}
wire w181;    //: /sn:0 {0}(809,2308)(809,2345)(828,2345)(828,2445){1}
wire w194;    //: /sn:0 {0}(682,2646)(682,2619)(681,2619)(681,2611){1}
wire w127;    //: /sn:0 {0}(965,1484)(965,1510)(981,1510)(981,1740){1}
wire w133;    //: /sn:0 {0}(707,2037)(707,1963)(673,1963)(673,1828)(694,1828)(694,1843)(709,1843)(709,1833){1}
//: {2}(709,1829)(709,1695){3}
//: {4}(707,1831)(694,1831)(694,1846){5}
wire w75;    //: /sn:0 {0}(512,973)(512,981)(515,981)(515,1004){1}
wire w204;    //: /sn:0 {0}(998,2875)(998,2774)(955,2774)(955,2636)(984,2636){1}
//: {2}(986,2634)(986,2541){3}
//: {4}(986,2638)(986,2650){5}
wire w276;    //: /sn:0 {0}(1101,3575)(1101,3549)(1285,3549)(1285,3405){1}
wire w209;    //: /sn:0 {0}(860,2677)(887,2677){1}
wire w215;    //: /sn:0 {0}(1052,2679)(1038,2679)(1038,2679)(1027,2679){1}
wire w156;    //: /sn:0 {0}(646,2377)(646,2348)(603,2348)(603,2224)(632,2224){1}
//: {2}(634,2222)(634,2055){3}
//: {4}(634,2226)(634,2240){5}
wire w41;    //: /sn:0 {0}(487,548)(487,556)(488,556)(488,575){1}
wire w36;    //: /sn:0 {0}(738,876)(738,709)(683,709)(683,567)(713,567){1}
//: {2}(715,565)(715,527)(744,527)(744,499){3}
//: {4}(715,569)(715,578){5}
wire w242;    //: /sn:0 {0}(994,3101)(964,3101){1}
wire w82;    //: /sn:0 {0}(501,1070)(501,1097)(526,1097)(526,1199){1}
wire w74;    //: /sn:0 {0}(391,1031)(370,1031)(370,1031)(362,1031){1}
wire w158;    //: /sn:0 {0}(968,1810)(968,1849){1}
wire w91;    //: /sn:0 {0}(760,1073)(760,1104)(786,1104)(786,1270){1}
wire w35;    //: /sn:0 {0}(651,850)(651,728)(602,728)(602,565)(630,565){1}
//: {2}(632,563)(632,507)(668,507)(668,474){3}
//: {4}(632,567)(632,577){5}
wire w101;    //: /sn:0 {0}(699,1653)(699,1538)(650,1538)(650,1397)(680,1397){1}
//: {2}(682,1395)(682,1300)(685,1300)(685,1289){3}
//: {4}(682,1399)(682,1415){5}
wire w163;    //: /sn:0 {0}(954,1915)(954,1949)(973,1949)(973,2111){1}
wire w265;    //: /sn:0 {0}(179,3412)(179,3374)(111,3374)(111,3307){1}
wire w22;    //: /sn:0 {0}(397,768)(397,747)(352,747)(352,563)(379,563){1}
//: {2}(381,561)(381,509)(422,509)(422,402){3}
//: {4}(381,565)(381,574){5}
wire w144;    //: /sn:0 {0}(576,2239)(576,2218)(577,2218)(577,2210){1}
wire w117;    //: /sn:0 {0}(890,1378)(890,1386)(891,1386)(891,1417){1}
wire w172;    //: /sn:0 {0}(660,2240)(660,2218)(659,2218)(659,2210){1}
wire w12;    //: /sn:0 {0}(419,133)(419,199){1}
wire w228;    //: /sn:0 {0}(827,3099)(807,3099)(807,3099)(802,3099){1}
wire w226;    //: /sn:0 {0}(1253,2719)(1253,2731)(1272,2731)(1272,2962){1}
wire w78;    //: /sn:0 {0}(593,973)(593,981)(595,981)(595,1005){1}
wire w200;    //: /sn:0 {0}(831,2816)(831,2767)(791,2767)(791,2637)(817,2637){1}
//: {2}(819,2635)(819,2487){3}
//: {4}(819,2639)(819,2648){5}
wire w257;    //: /sn:0 {0}(331,741)(331,702)(312,702)(312,639){1}
wire w27;    //: /sn:0 {0}(688,231)(674,231)(674,231)(668,231){1}
wire w86;    //: /sn:0 {0}(734,1035)(708,1035)(708,1035)(697,1035){1}
wire w138;    //: /sn:0 {0}(459,1924)(459,1909){1}
wire w246;    //: /sn:0 {0}(1114,3074)(1114,3039)(1113,3039)(1113,3031){1}
wire w80;    //: /sn:0 {0}(555,1033)(545,1033)(545,1033)(530,1033){1}
wire w29;    //: /sn:0 {0}(639,268)(639,298)(677,298)(677,432){1}
wire w231;    //: /sn:0 {0}(935,3261)(935,3186)(892,3186)(892,3057)(921,3057){1}
//: {2}(923,3055)(923,2887){3}
//: {4}(923,3059)(923,3072){5}
wire w264;    //: /sn:0 {0}(189,3412)(189,3324)(163,3324)(163,3307){1}
wire w42;    //: /sn:0 {0}(300,573)(300,559){1}
//: {2}(300,555)(300,503)(334,503)(334,380){3}
//: {4}(298,557)(272,557)(272,722)(312,722)(312,741){5}
wire w147;    //: /sn:0 {0}(624,1911)(624,1942)(643,1942)(643,2013){1}
wire w277;    //: /sn:0 {0}(1111,3575)(1111,3556)(1375,3556)(1375,3429){1}
wire w247;    //: /sn:0 {0}(1020,3139)(1020,3169)(1039,3169)(1039,3290){1}
wire w112;    //: /sn:0 {0}(516,1479)(516,1510)(541,1510)(541,1588){1}
wire w60;    //: /sn:0 {0}(821,645)(821,671)(831,671)(831,903){1}
wire w46;    //: /sn:0 {0}(534,604)(504,604)(504,604)(503,604){1}
wire w175;    //: /sn:0 {0}(646,2306)(646,2337)(665,2337)(665,2377){1}
wire w15;    //: /sn:0 {0}(458,228)(434,228){1}
wire w109;    //: /sn:0 {0}(435,1478)(435,1499)(454,1499)(454,1559){1}
wire w129;    //: /sn:0 {0}(515,1872)(495,1872)(495,1872)(488,1872){1}
wire w114;    //: /sn:0 {0}(796,1378)(796,1386)(799,1386)(799,1416){1}
wire w97;    //: /sn:0 {0}(62,3265)(62,3232)(85,3232)(85,718){1}
//: {2}(87,716)(99,716)(99,717)(144,717)(144,763){3}
//: {4}(146,765)(297,765){5}
//: {6}(144,767)(144,790){7}
//: {8}(146,792)(382,792){9}
//: {10}(144,794)(144,818){11}
//: {12}(146,820)(465,820){13}
//: {14}(144,822)(144,844){15}
//: {16}(146,846)(550,846){17}
//: {18}(144,848)(144,872){19}
//: {20}(146,874)(636,874){21}
//: {22}(144,876)(144,898){23}
//: {24}(146,900)(723,900){25}
//: {26}(144,902)(144,927)(797,927){27}
//: {28}(85,714)(85,600)(201,600){29}
wire w229;    //: /sn:0 {0}(773,3209)(773,3179)(728,3179)(728,3054)(759,3054){1}
//: {2}(761,3052)(761,2809){3}
//: {4}(761,3056)(761,3070){5}
wire w267;    //: /sn:0 {0}(159,3412)(159,3392)(9,3392)(9,3307){1}
wire w261;    //: /sn:0 {0}(219,3412)(219,3385)(331,3385)(331,3308){1}
wire w64;    //: /sn:0 {0}(367,1378)(367,1386)(369,1386)(369,1411){1}
wire w245;    //: /sn:0 {0}(1074,3102)(1049,3102){1}
wire w259;    //: /sn:0 {0}(1365,3143)(1365,3171)(1384,3171)(1384,3387){1}
wire w63;    //: /sn:0 {0}(236,1001)(236,936)(322,936)(322,783){1}
wire w159;    //: /sn:0 {0}(869,1914)(869,1947)(888,1947)(888,2088){1}
wire w76;    //: /sn:0 {0}(333,1068)(333,1084)(352,1084)(352,1141){1}
wire w21;    //: /sn:0 {0}(515,384)(515,288)(484,288)(484,266){1}
wire w236;    //: /sn:0 {0}(1350,3411)(633,3411)(633,3389){1}
//: {2}(635,3387)(1260,3387){3}
//: {4}(633,3385)(633,3367){5}
//: {6}(635,3365)(1170,3365){7}
//: {8}(633,3363)(633,3345){9}
//: {10}(635,3343)(1085,3343){11}
//: {12}(633,3341)(633,3316){13}
//: {14}(635,3314)(1005,3314){15}
//: {16}(633,3312)(633,3287){17}
//: {18}(635,3285)(920,3285){19}
//: {20}(633,3283)(633,3260){21}
//: {22}(635,3258)(838,3258){23}
//: {24}(633,3256)(633,3235){25}
//: {26}(635,3233)(758,3233){27}
//: {28}(633,3231)(633,3100){29}
//: {30}(635,3098)(747,3098){31}
//: {32}(631,3098)(385,3098)(385,3266){33}
wire w170;    //: /sn:0 {0}(276,3266)(276,3251)(246,3251)(246,2401){1}
//: {2}(248,2399)(256,2399)(256,2401)(506,2401){3}
//: {4}(510,2401)(631,2401){5}
//: {6}(508,2403)(508,2435){7}
//: {8}(510,2437)(714,2437){9}
//: {10}(508,2439)(508,2467){11}
//: {12}(510,2469)(794,2469){13}
//: {14}(508,2471)(508,2496){15}
//: {16}(510,2498)(876,2498){17}
//: {18}(508,2500)(508,2521){19}
//: {20}(510,2523)(961,2523){21}
//: {22}(508,2525)(508,2549){23}
//: {24}(510,2551)(1041,2551){25}
//: {26}(508,2553)(508,2575)(1126,2575){27}
//: {28}(246,2397)(246,2267)(536,2267){29}
wire w199;    //: /sn:0 {0}(1163,2930)(1163,2784)(1122,2784)(1122,2641)(1149,2641){1}
//: {2}(1151,2639)(1151,2593){3}
//: {4}(1151,2643)(1151,2652){5}
wire w100;    //: /sn:0 {0}(610,1624)(610,1514)(559,1514)(559,1393)(591,1393){1}
//: {2}(593,1391)(593,1277)(599,1277)(599,1266){3}
//: {4}(593,1395)(593,1414){5}
wire w230;    //: /sn:0 {0}(853,3234)(853,3180)(812,3180)(812,3055)(839,3055){1}
//: {2}(841,3053)(841,2858){3}
//: {4}(841,3057)(841,3071){5}
wire w249;    //: /sn:0 {0}(1199,3075)(1199,3031){1}
wire w24;    //: /sn:0 {0}(652,133)(652,141)(653,141)(653,202){1}
wire w251;    //: /sn:0 {0}(1249,3104)(1214,3104){1}
wire w260;    //: /sn:0 {0}(386,3308)(386,3394)(229,3394)(229,3412){1}
wire w256;    //: /sn:0 {0}(1275,3142)(1275,3165)(1294,3165)(1294,3363){1}
wire w1;    //: /sn:0 {0}(242,548)(242,556)(241,556)(241,572){1}
wire w161;    //: /sn:0 {0}(1008,1878)(996,1878)(996,1878)(983,1878){1}
wire w140;    //: /sn:0 {0}(1141,2551)(1141,2398)(1099,2398)(1099,2226)(1127,2226){1}
//: {2}(1129,2224)(1129,1227)(1357,1227){3}
//: {4}(1129,2228)(1129,2246){5}
wire w196;    //: /sn:0 {0}(656,2646)(656,2436)(656,2436)(656,2419){1}
wire w221;    //: /sn:0 {0}(1227,2681)(1192,2681){1}
wire w235;    //: /sn:0 {0}(1275,3363)(1275,3205)(1228,3205)(1228,3060)(1261,3060){1}
//: {2}(1263,3058)(1263,3004){3}
//: {4}(1263,3062)(1263,3076){5}
wire w241;    //: /sn:0 {0}(853,3137)(853,3167)(872,3167)(872,3234){1}
wire w154;    //: /sn:0 {0}(882,1810)(882,1818)(883,1818)(883,1848){1}
wire w205;    //: /sn:0 {0}(765,2647)(765,2619)(764,2619)(764,2611){1}
wire w253;    //: /sn:0 {0}(1185,3141)(1185,3173)(1204,3173)(1204,3341){1}
wire w116;    //: /sn:0 {0}(759,1444)(723,1444){1}
wire w98;    //: /sn:0 {0}(435,1559)(435,1509)(393,1509)(393,1400)(421,1400){1}
//: {2}(423,1398)(423,1223)(428,1223)(428,1210){3}
//: {4}(423,1402)(423,1412){5}
wire w227;    //: /sn:0 {0}(787,3070)(787,3039)(786,3039)(786,3031){1}
wire w18;    //: /sn:0 {0}(541,1984)(541,1936)(503,1936)(503,1829)(527,1829){1}
//: {2}(531,1829)(532,1829)(532,1630){3}
//: {4}(529,1831)(529,1844){5}
wire w118;    //: /sn:0 {0}(694,1481)(694,1509)(718,1509)(718,1653){1}
wire w212;    //: /sn:0 {0}(972,2678)(942,2678){1}
wire w243;    //: /sn:0 {0}(1034,3073)(1034,3039)(1033,3039)(1033,3031){1}
wire w164;    //: /sn:0 {0}(1034,2135)(1034,2012)(993,2012)(993,1834)(1020,1834){1}
//: {2}(1022,1832)(1022,740)(1357,740){3}
//: {4}(1022,1836)(1022,1850){5}
wire w68;    //: /sn:0 {0}(447,1378)(447,1386)(449,1386)(449,1412){1}
wire w198;    //: /sn:0 {0}(751,2767)(751,2751)(712,2751)(712,2631)(737,2631){1}
//: {2}(739,2629)(739,2455){3}
//: {4}(739,2633)(739,2647){5}
wire w123;    //: /sn:0 {0}(962,1740)(962,1529)(923,1529)(923,1405)(951,1405){1}
//: {2}(953,1403)(953,584)(1357,584){3}
//: {4}(953,1407)(953,1418){5}
wire w62;    //: /sn:0 {0}(307,1030)(289,1030)(289,1030)(277,1030){1}
wire w85;    //: /sn:0 {0}(581,1071)(581,1101)(608,1101)(608,1224){1}
wire w185;    //: /sn:0 {0}(1030,2273)(1015,2273)(1015,2273)(1005,2273){1}
wire w137;    //: /sn:0 {0}(217,3266)(217,3245)(194,3245)(194,2009){1}
//: {2}(196,2007)(204,2007)(204,2008)(252,2008){3}
//: {4}(256,2008)(526,2008){5}
//: {6}(254,2010)(254,2035){7}
//: {8}(256,2037)(609,2037){9}
//: {10}(254,2039)(254,2059){11}
//: {12}(256,2061)(692,2061){13}
//: {14}(254,2063)(254,2084){15}
//: {16}(256,2086)(772,2086){17}
//: {18}(254,2088)(254,2110){19}
//: {20}(256,2112)(854,2112){21}
//: {22}(254,2114)(254,2133){23}
//: {24}(256,2135)(939,2135){25}
//: {26}(254,2137)(254,2159)(1019,2159){27}
//: {28}(194,2005)(194,1871)(433,1871){29}
wire w11;    //: /sn:0 {0}(379,227)(363,227)(363,227)(354,227){1}
wire w197;    //: /sn:0 {0}(1078,2903)(1078,2773)(1037,2773)(1037,2630)(1064,2630){1}
//: {2}(1066,2628)(1066,2569){3}
//: {4}(1066,2632)(1066,2651){5}
wire w150;    //: /sn:0 {0}(784,1810)(784,1818)(801,1818)(801,1847){1}
wire w70;    //: /sn:0 {0}(767,1270)(767,1144)(712,1144)(712,995)(746,995){1}
//: {2}(748,993)(748,958)(822,958)(822,945){3}
//: {4}(748,997)(748,1007){5}
wire w110;    //: /sn:0 {0}(579,1442)(545,1442){1}
wire w189;    //: /sn:0 {0}(1155,2246)(1155,2218)(1154,2218)(1154,2210){1}
wire w193;    //: /sn:0 {0}(1141,2312)(1141,2337)(1160,2337)(1160,2551){1}
wire w206;    //: /sn:0 {0}(805,2676)(792,2676)(792,2676)(780,2676){1}
wire w13;    //: /sn:0 {0}(325,264)(325,291)(343,291)(343,338){1}
wire w88;    //: /sn:0 {0}(668,1072)(668,1097)(694,1097)(694,1247){1}
wire w5;    //: /sn:0 {0}(254,133)(254,141)(256,141)(256,197){1}
wire w48;    //: /sn:0 {0}(499,796)(499,666)(474,666)(474,641){1}
wire w208;    //: /sn:0 {0}(751,2713)(751,2736)(770,2736)(770,2767){1}
wire w131;    //: /sn:0 {0}(624,2013)(624,1967)(582,1967)(582,1846)(620,1846)(620,1834){1}
//: {2}(620,1830)(620,1666){3}
//: {4}(618,1832)(612,1832)(612,1845){5}
wire w47;    //: /sn:0 {0}(658,548)(658,577){1}
wire w26;    //: /sn:0 {0}(480,796)(480,695)(433,695)(433,563)(460,563){1}
//: {2}(462,561)(462,513)(506,513)(506,426){3}
//: {4}(462,565)(462,575){5}
//: enddecls

  FS g8 (.A(w31), .B(w24), .Bin(w27), .Bout(w23), .D(w29));   //: @(614, 203) /sz:(53, 64) /sn:0 /p:[ Ti0>43 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FS g165 (.A(w18), .B(w139), .Bin(w141), .Bout(w129), .D(w132));   //: @(516, 1845) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w44 = B[3]; //: TAP g55 @(573,542) /sn:0 /R:1 /w:[ 0 26 25 ] /ss:1
  MUX2 g37 (.in0(w29), .in1(w31), .c(w3), .out(w35));   //: @(644, 433) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>3 Bo0<3 ]
  assign w0 = B[7]; //: TAP g13 @(169,127) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: GROUND g140 (w126) @(1009,1421) /sn:0 /R:2 /w:[ 0 ]
  assign w68 = B[6]; //: TAP g139 @(447,1372) /sn:0 /R:1 /w:[ 0 68 67 ] /ss:1
  //: OUT g310 (D) @(235,3436) /sn:0 /w:[ 0 ]
  MUX2 g111 (.in0(w85), .in1(w67), .c(w71), .out(w100));   //: @(575, 1225) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>17 Bo0<3 ]
  MUX2 g314 (.in1(w230), .in0(w241), .c(w236), .out(w271));   //: @(839, 3235) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>23 Bo0<1 ]
  assign w150 = B[3]; //: TAP g176 @(784,1804) /sn:0 /R:1 /w:[ 0 81 82 ] /ss:1
  assign w189 = B[0]; //: TAP g218 @(1154,2204) /sn:0 /R:1 /w:[ 1 107 108 ] /ss:1
  //: IN g1 (B) @(56,129) /sn:0 /w:[ 0 ]
  //: joint g328 (w231) @(923, 3057) /w:[ -1 2 1 4 ]
  //: joint g277 (w201) @(550, 2927) /w:[ 20 19 -1 22 ]
  assign w30 = A[7]; //: TAP g11 @(700,80) /sn:0 /R:1 /w:[ 3 1 2 ] /ss:1
  FS g130 (.A(w102), .B(w114), .Bin(w119), .Bout(w116), .D(w121));   //: @(760, 1417) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  INV1 g306 (.in(w71), .out(w265));   //: @(91, 3266) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  //: joint g266 (w201) @(550, 2791) /w:[ 4 -1 3 6 ]
  FS g50 (.A(w36), .B(w50), .Bin(w55), .Bout(w52), .D(w57));   //: @(702, 579) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  FS g254 (.B(w216), .A(w197), .Bin(w218), .Bout(w215), .D(w220));   //: @(1053, 2652) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g223 (w140) @(1129, 2226) /w:[ -1 2 1 4 ]
  //: joint g113 (w67) @(569, 994) /w:[ -1 2 1 4 ]
  assign w24 = B[1]; //: TAP g19 @(652,127) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  FS g132 (.A(w123), .B(w120), .Bin(w126), .Bout(w122), .D(w127));   //: @(940, 1419) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g197 (.in1(w136), .in0(w163), .c(w137), .out(w168));   //: @(940, 2112) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>25 Bo0<3 ]
  //: joint g330 (w230) @(841, 3055) /w:[ -1 2 1 4 ]
  //: joint g150 (w100) @(593, 1393) /w:[ -1 2 1 4 ]
  //: joint g146 (w104) @(157, 1583) /w:[ 2 28 -1 1 ]
  //: joint g38 (w31) @(393, 189) /w:[ -1 29 30 32 ]
  INV1 g307 (.in(w97), .out(w266));   //: @(43, 3266) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  //: joint g115 (w71) @(142, 1248) /w:[ 16 15 -1 18 ]
  //: joint g75 (w97) @(144, 820) /w:[ 12 11 -1 14 ]
  //: joint g227 (w168) @(964, 2226) /w:[ -1 2 1 4 ]
  MUX2 g31 (.in0(w17), .in1(w31), .c(w3), .out(w22));   //: @(398, 361) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>31 Li0>15 Bo0<3 ]
  //: GROUND g20 (w31) @(107,174) /sn:0 /R:3 /w:[ 21 ]
  assign w114 = B[2]; //: TAP g135 @(796,1372) /sn:0 /R:1 /w:[ 0 60 59 ] /ss:1
  MUX2 g160 (.in0(w127), .in1(w123), .c(w104), .out(w136));   //: @(948, 1741) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>27 Bo0<3 ]
  FS g169 (.A(w135), .B(w154), .Bin(w157), .Bout(w153), .D(w159));   //: @(844, 1849) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FS g124 (.A(w95), .B(w64), .Bin(w92), .Bout(w104), .D(w105));   //: @(330, 1412) /sz:(53, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<29 Bo0<1 ]
  MUX2 g230 (.in1(w168), .in0(w187), .c(w170), .out(w204));   //: @(962, 2500) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>21 Bo0<3 ]
  //: joint g68 (w97) @(144, 765) /w:[ 4 3 -1 6 ]
  //: joint g39 (w3) @(206, 433) /w:[ 6 8 -1 5 ]
  assign w227 = B[7]; //: TAP g284 @(786,3025) /sn:0 /R:1 /w:[ 1 131 132 ] /ss:1
  //: joint g195 (w135) @(857, 1831) /w:[ -1 2 1 4 ]
  //: joint g107 (w71) @(142, 1165) /w:[ 4 -1 3 6 ]
  assign w53 = B[0]; //: TAP g52 @(807,542) /sn:0 /R:1 /w:[ 0 20 19 ] /ss:1
  assign w162 = B[0]; //: TAP g179 @(1049,1804) /sn:0 /R:1 /w:[ 0 87 88 ] /ss:1
  FS g205 (.B(w172), .A(w156), .Bin(w173), .Bout(w148), .D(w175));   //: @(621, 2241) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g231 (w165) @(797, 2231) /w:[ -1 2 1 4 ]
  //: joint g201 (w164) @(1022, 1834) /w:[ -1 2 1 4 ]
  FS g297 (.B(w255), .A(w224), .Bin(w258), .Bout(w254), .D(w259));   //: @(1340, 3078) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g221 (.in1(w198), .in0(w208), .c(w201), .out(w229));   //: @(737, 2768) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>5 Bo0<3 ]
  //: joint g321 (w236) @(633, 3285) /w:[ 18 20 -1 17 ]
  MUX2 g320 (.in1(w232), .in0(w247), .c(w236), .out(w273));   //: @(1006, 3291) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>15 Bo0<1 ]
  assign w5 = B[6]; //: TAP g14 @(254,127) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  FS g47 (.A(w26), .B(w41), .Bin(w46), .Bout(w43), .D(w48));   //: @(449, 576) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  FS g44 (.A(w14), .B(w1), .Bin(w10), .Bout(w97), .D(w38));   //: @(202, 573) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<29 Bo0<1 ]
  //: joint g84 (w56) @(817, 564) /w:[ 2 1 4 -1 ]
  MUX2 g105 (.in0(w79), .in1(w66), .c(w71), .out(w98));   //: @(404, 1169) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>9 Bo0<3 ]
  assign w205 = B[6]; //: TAP g247 @(764,2605) /sn:0 /R:1 /w:[ 1 115 116 ] /ss:1
  //: joint g23 (w31) @(313, 174) /w:[ 11 12 14 26 ]
  //: joint g236 (w170) @(508, 2498) /w:[ 16 15 -1 18 ]
  //: joint g116 (w96) @(489, 989) /w:[ -1 2 1 4 ]
  MUX2 g311 (.in1(w229), .in0(w237), .c(w236), .out(w270));   //: @(759, 3210) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>27 Bo0<1 ]
  FS g93 (.A(w96), .B(w75), .Bin(w80), .Bout(w77), .D(w82));   //: @(476, 1005) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w47 = B[2]; //: TAP g54 @(658,542) /sn:0 /R:1 /w:[ 0 24 23 ] /ss:1
  MUX2 g40 (.in0(w33), .in1(w30), .c(w3), .out(w36));   //: @(720, 458) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Bo0<3 ]
  assign w207 = B[5]; //: TAP g249 @(844,2605) /sn:0 /R:1 /w:[ 1 117 118 ] /ss:1
  //: joint g337 (w31) @(627, 182) /w:[ -1 2 1 42 ]
  FS g46 (.A(w22), .B(w39), .Bin(w43), .Bout(w40), .D(w45));   //: @(368, 575) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g26 (w31) @(550, 174) /w:[ 3 4 6 40 ]
  //: IN g0 (A) @(56,82) /sn:0 /w:[ 0 ]
  FS g167 (.A(w133), .B(w146), .Bin(w149), .Bout(w145), .D(w151));   //: @(681, 1847) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g316 (w235) @(1263, 3060) /w:[ -1 2 1 4 ]
  //: joint g278 (w199) @(1151, 2641) /w:[ -1 2 1 4 ]
  MUX2 g228 (.in1(w166), .in0(w184), .c(w170), .out(w202));   //: @(877, 2475) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>17 Bo0<3 ]
  assign w111 = B[3]; //: TAP g136 @(706,1372) /sn:0 /R:1 /w:[ 0 62 61 ] /ss:1
  MUX2 g224 (.in1(w160), .in0(w178), .c(w170), .out(w198));   //: @(715, 2414) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>9 Bo0<3 ]
  //: joint g233 (w170) @(508, 2401) /w:[ 4 -1 3 6 ]
  assign w139 = B[6]; //: TAP g173 @(554,1804) /sn:0 /R:1 /w:[ 0 75 76 ] /ss:1
  //: joint g190 (w137) @(254, 2037) /w:[ 8 7 -1 10 ]
  //: GROUND g61 (w37) @(894,1015) /sn:0 /R:2 /w:[ 0 ]
  //: joint g331 (w236) @(633, 3365) /w:[ 6 8 -1 5 ]
  //: joint g86 (B) @(115, 969) /w:[ 36 35 -1 150 ]
  //: joint g34 (w3) @(206, 384) /w:[ 14 16 -1 13 ]
  FS g3 (.A(w31), .B(w5), .Bin(w7), .Bout(w2), .D(w9));   //: @(217, 198) /sz:(53, 64) /sn:0 /p:[ Ti0>25 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w140 = A[2]; //: TAP g220 @(1360,1227) /sn:0 /R:2 /w:[ 3 12 11 ] /ss:0
  MUX2 g267 (.in1(w202), .in0(w214), .c(w201), .out(w231));   //: @(899, 2846) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>13 Bo0<3 ]
  assign w191 = A[1]; //: TAP g261 @(1360,2385) /sn:0 /R:2 /w:[ 3 14 13 ] /ss:0
  //: joint g110 (w71) @(142, 1192) /w:[ 8 7 -1 10 ]
  assign w90 = A[5]; //: TAP g65 @(1360,360) /sn:0 /R:2 /w:[ 3 6 5 ] /ss:0
  FS g250 (.B(w210), .A(w202), .Bin(w212), .Bout(w209), .D(w214));   //: @(888, 2650) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<1 Bo0<0 ]
  assign w1 = B[7]; //: TAP g59 @(242,542) /sn:0 /R:1 /w:[ 0 34 33 ] /ss:1
  //: joint g147 (w104) @(363, 1583) /w:[ 4 -1 3 6 ]
  //: joint g156 (w104) @(363, 1677) /w:[ 16 15 -1 18 ]
  //: joint g325 (w232) @(1008, 3060) /w:[ -1 2 1 4 ]
  //: joint g153 (w104) @(363, 1648) /w:[ 12 11 -1 14 ]
  assign w81 = B[2]; //: TAP g98 @(681,967) /sn:0 /R:1 /w:[ 0 47 48 ] /ss:1
  MUX2 g317 (.in1(w231), .in0(w244), .c(w236), .out(w272));   //: @(921, 3262) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>19 Bo0<1 ]
  INV1 g304 (.in(w137), .out(w263));   //: @(198, 3267) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  assign w78 = B[3]; //: TAP g96 @(593,967) /sn:0 /R:1 /w:[ 0 45 46 ] /ss:1
  assign w12 = B[4]; //: TAP g16 @(419,127) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: joint g183 (w18) @(529, 1829) /w:[ 2 -1 1 4 ]
  //: joint g122 (w65) @(321, 988) /w:[ -1 2 1 4 ]
  //: joint g280 (w191) @(1241, 2641) /w:[ -1 2 1 4 ]
  FS g87 (.A(w63), .B(w58), .Bin(w62), .Bout(w71), .D(w72));   //: @(223, 1002) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<29 Bo0<1 ]
  //: joint g78 (w97) @(144, 846) /w:[ 16 15 -1 18 ]
  FS g129 (.A(w101), .B(w111), .Bin(w116), .Bout(w113), .D(w118));   //: @(669, 1416) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FS g171 (.A(w164), .B(w162), .Bin(w128), .Bout(w161), .D(w167));   //: @(1009, 1851) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FS g258 (.B(w222), .A(w191), .Bin(w225), .Bout(w221), .D(w226));   //: @(1228, 2654) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g143 (w98) @(423, 1400) /w:[ -1 2 1 4 ]
  //: joint g69 (w22) @(381, 563) /w:[ -1 2 1 4 ]
  INV1 g305 (.in(w104), .out(w264));   //: @(143, 3266) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  FS g244 (.B(w194), .A(w196), .Bin(w195), .Bout(w201), .D(w203));   //: @(643, 2647) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<29 Bo0<0 ]
  //: joint g119 (w71) @(142, 1271) /w:[ 20 19 -1 22 ]
  assign w194 = B[7]; //: TAP g245 @(681,2605) /sn:0 /R:1 /w:[ 1 113 114 ] /ss:1
  assign w8 = B[5]; //: TAP g15 @(335,127) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g162 (w123) @(953, 1405) /w:[ -1 2 1 4 ]
  INV1 g308 (.in(w3), .out(w267));   //: @(-11, 3266) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>29 Bo0<1 ]
  //: joint g322 (w233) @(1088, 3059) /w:[ -1 2 1 4 ]
  FS g131 (.A(w103), .B(w117), .Bin(w122), .Bout(w119), .D(w124));   //: @(852, 1418) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g67 (.in0(w45), .in1(w22), .c(w97), .out(w65));   //: @(383, 769) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>9 Bo0<3 ]
  FS g127 (.A(w99), .B(w106), .Bin(w110), .Bout(w107), .D(w112));   //: @(491, 1414) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FS g293 (.B(w249), .A(w234), .Bin(w251), .Bout(w248), .D(w253));   //: @(1160, 3076) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<1 Bo0<0 ]
  //: joint g43 (B) @(826, 544) /w:[ -1 17 18 152 ]
  //: joint g315 (w236) @(633, 3233) /w:[ 26 28 -1 25 ]
  //: joint g62 (w97) @(85, 716) /w:[ 2 28 -1 1 ]
  assign w58 = B[7]; //: TAP g88 @(260,967) /sn:0 /R:1 /w:[ 0 37 38 ] /ss:1
  //: joint g104 (w71) @(112, 1165) /w:[ 2 28 -1 1 ]
  assign w106 = B[5]; //: TAP g138 @(530,1372) /sn:0 /R:1 /w:[ 0 66 65 ] /ss:1
  assign w87 = B[0]; //: TAP g63 @(861,967) /sn:0 /R:1 /w:[ 0 51 52 ] /ss:1
  MUX2 g188 (.in1(w133), .in0(w151), .c(w137), .out(w160));   //: @(693, 2038) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>13 Bo0<3 ]
  assign w219 = B[1]; //: TAP g257 @(1176,2605) /sn:0 /R:1 /w:[ 1 125 126 ] /ss:1
  //: joint g109 (w69) @(656, 994) /w:[ -1 2 1 4 ]
  assign w146 = B[4]; //: TAP g175 @(720,1804) /sn:0 /R:1 /w:[ 0 79 80 ] /ss:1
  //: joint g234 (w170) @(508, 2437) /w:[ 8 7 -1 10 ]
  FS g285 (.B(w238), .A(w230), .Bin(w239), .Bout(w228), .D(w241));   //: @(828, 3072) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g264 (.in1(w200), .in0(w211), .c(w201), .out(w230));   //: @(817, 2817) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>9 Bo0<3 ]
  assign w120 = B[0]; //: TAP g133 @(978,1372) /sn:0 /R:1 /w:[ 0 56 55 ] /ss:1
  FS g5 (.A(w31), .B(w12), .Bin(w15), .Bout(w11), .D(w17));   //: @(380, 200) /sz:(53, 64) /sn:0 /p:[ Ti0>33 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w41 = B[4]; //: TAP g56 @(487,542) /sn:0 /R:1 /w:[ 0 28 27 ] /ss:1
  FS g95 (.A(w67), .B(w78), .Bin(w83), .Bout(w80), .D(w85));   //: @(556, 1006) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g24 (w31) @(395, 174) /w:[ 9 -1 10 28 ]
  //: GROUND g85 (w59) @(880,589) /sn:0 /R:2 /w:[ 0 ]
  assign w73 = B[5]; //: TAP g92 @(431,967) /sn:0 /R:1 /w:[ 0 41 42 ] /ss:1
  //: joint g333 (w229) @(761, 3054) /w:[ -1 2 1 4 ]
  //: joint g313 (w236) @(633, 3098) /w:[ 30 -1 32 29 ]
  assign w56 = A[6]; //: TAP g60 @(929,80) /sn:0 /R:1 /w:[ 3 3 4 ] /ss:1
  FS g101 (.A(w90), .B(w87), .Bin(w37), .Bout(w89), .D(w94));   //: @(823, 1008) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w177 = B[4]; //: TAP g210 @(821,2204) /sn:0 /R:1 /w:[ 1 99 100 ] /ss:1
  assign w183 = B[2]; //: TAP g214 @(989,2204) /sn:0 /R:1 /w:[ 1 103 104 ] /ss:1
  MUX2 g332 (.in1(w224), .in0(w259), .c(w236), .out(w277));   //: @(1351, 3388) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>0 Bo0<1 ]
  INV1 g303 (.in(w170), .out(w262));   //: @(255, 3267) /sz:(41, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  FS g170 (.A(w136), .B(w158), .Bin(w161), .Bout(w157), .D(w163));   //: @(929, 1850) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g35 (.in0(w25), .in1(w31), .c(w3), .out(w34));   //: @(564, 410) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>5 Li0>7 Bo0<3 ]
  FS g126 (.A(w98), .B(w68), .Bin(w107), .Bout(w92), .D(w109));   //: @(410, 1413) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g185 (.in1(w131), .in0(w147), .c(w137), .out(w156));   //: @(610, 2014) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>9 Bo0<3 ]
  assign w144 = B[7]; //: TAP g204 @(577,2204) /sn:0 /R:1 /w:[ 1 93 94 ] /ss:1
  assign w210 = B[4]; //: TAP g251 @(926,2605) /sn:0 /R:1 /w:[ 1 119 120 ] /ss:1
  //: joint g66 (w42) @(300, 557) /w:[ -1 2 4 1 ]
  FS g97 (.A(w69), .B(w81), .Bin(w86), .Bout(w83), .D(w88));   //: @(643, 1007) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g120 (.in0(w94), .in1(w90), .c(w71), .out(w103));   //: @(836, 1296) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>27 Bo0<3 ]
  //: joint g184 (w137) @(194, 2007) /w:[ 2 28 -1 1 ]
  //: joint g235 (w170) @(508, 2469) /w:[ 12 11 -1 14 ]
  //: GROUND g260 (w225) @(1304,2655) /sn:0 /R:2 /w:[ 0 ]
  assign w28 = B[0]; //: TAP g12 @(728,127) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  assign w20 = B[2]; //: TAP g18 @(577,127) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  MUX2 g226 (.in1(w165), .in0(w181), .c(w170), .out(w200));   //: @(795, 2446) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>13 Bo0<3 ]
  //: joint g239 (w160) @(717, 2228) /w:[ -1 2 1 4 ]
  FS g283 (.B(w227), .A(w229), .Bin(w228), .Bout(w236), .D(w237));   //: @(748, 3071) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<31 Bo0<0 ]
  MUX2 g108 (.in0(w82), .in1(w96), .c(w71), .out(w99));   //: @(493, 1200) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>13 Bo0<3 ]
  MUX2 g191 (.in1(w134), .in0(w155), .c(w137), .out(w165));   //: @(773, 2063) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>17 Bo0<3 ]
  //: GROUND g219 (w192) @(1186,2247) /sn:0 /R:2 /w:[ 0 ]
  //: OUT g336 (R) @(1109,3623) /sn:0 /w:[ 0 ]
  MUX2 g326 (.in1(w234), .in0(w253), .c(w236), .out(w275));   //: @(1171, 3342) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>7 Bo0<1 ]
  assign w117 = B[1]; //: TAP g134 @(890,1372) /sn:0 /R:1 /w:[ 0 58 57 ] /ss:1
  //: joint g242 (w170) @(508, 2551) /w:[ 24 23 -1 26 ]
  //: joint g281 (w201) @(550, 2954) /w:[ 24 23 -1 26 ]
  FS g4 (.A(w31), .B(w8), .Bin(w11), .Bout(w7), .D(w13));   //: @(300, 199) /sz:(53, 64) /sn:0 /p:[ Ti0>27 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g154 (.in0(w121), .in1(w102), .c(w104), .out(w134));   //: @(774, 1683) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>21 Bo0<3 ]
  MUX2 g237 (.in1(w169), .in0(w190), .c(w170), .out(w197));   //: @(1042, 2528) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>25 Bo0<3 ]
  //: joint g186 (w131) @(620, 1832) /w:[ -1 2 4 1 ]
  assign w6 = B[6]; //: TAP g58 @(326,542) /sn:0 /R:1 /w:[ 0 32 31 ] /ss:1
  //: joint g112 (w71) @(142, 1223) /w:[ 12 11 -1 14 ]
  //: joint g268 (w201) @(550, 2840) /w:[ 8 7 -1 10 ]
  MUX2 g76 (.in0(w54), .in1(w35), .c(w97), .out(w67));   //: @(637, 851) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>21 Bo0<3 ]
  FS g211 (.B(w180), .A(w166), .Bin(w182), .Bout(w179), .D(w184));   //: @(866, 2244) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g319 (w234) @(1173, 3061) /w:[ -1 2 1 4 ]
  //: joint g324 (w236) @(633, 3314) /w:[ 14 16 -1 13 ]
  assign w246 = B[3]; //: TAP g292 @(1113,3025) /sn:0 /R:1 /w:[ 1 139 140 ] /ss:1
  MUX2 g157 (.in0(w124), .in1(w103), .c(w104), .out(w135));   //: @(869, 1713) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>25 Bo0<3 ]
  //: joint g163 (B) @(279, 1806) /w:[ 72 71 -1 90 ]
  //: joint g238 (w170) @(508, 2523) /w:[ 20 19 -1 22 ]
  assign R = {w270, w271, w272, w273, w274, w275, w276, w277}; //: CONCAT g335  @(1076,3580) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g263 (w201) @(325, 2790) /w:[ 2 28 -1 1 ]
  assign w222 = B[0]; //: TAP g259 @(1266,2605) /sn:0 /R:1 /w:[ 1 127 128 ] /ss:1
  MUX2 g64 (.in0(w257), .in1(w42), .c(w97), .out(w63));   //: @(298, 742) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>5 Li0>5 Bo0<1 ]
  FS g166 (.A(w131), .B(w142), .Bin(w145), .Bout(w141), .D(w147));   //: @(599, 1846) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g241 (w156) @(634, 2224) /w:[ -1 2 1 4 ]
  //: joint g334 (w236) @(633, 3387) /w:[ 2 4 -1 1 ]
  assign w249 = B[2]; //: TAP g294 @(1199,3025) /sn:0 /R:1 /w:[ 1 141 142 ] /ss:1
  //: joint g274 (w201) @(550, 2899) /w:[ 16 15 -1 18 ]
  //: joint g121 (w71) @(142, 1294) /w:[ 24 23 -1 26 ]
  assign w172 = B[6]; //: TAP g206 @(659,2204) /sn:0 /R:1 /w:[ 1 95 96 ] /ss:1
  //: joint g28 (w3) @(42, 333) /w:[ 25 26 -1 28 ]
  //: joint g225 (w169) @(1044, 2230) /w:[ -1 2 1 4 ]
  //: joint g265 (w200) @(819, 2637) /w:[ -1 2 1 4 ]
  //: joint g272 (w201) @(550, 2869) /w:[ 12 11 -1 14 ]
  FS g6 (.A(w31), .B(w16), .Bin(w19), .Bout(w15), .D(w21));   //: @(459, 201) /sz:(53, 64) /sn:0 /p:[ Ti0>39 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  assign w154 = B[2]; //: TAP g177 @(882,1804) /sn:0 /R:1 /w:[ 0 83 84 ] /ss:1
  //: joint g192 (w137) @(254, 2061) /w:[ 12 11 -1 14 ]
  assign w174 = B[5]; //: TAP g208 @(743,2204) /sn:0 /R:1 /w:[ 1 97 98 ] /ss:1
  assign w50 = B[1]; //: TAP g53 @(738,542) /sn:0 /R:1 /w:[ 0 22 21 ] /ss:1
  FS g7 (.A(w31), .B(w20), .Bin(w23), .Bout(w19), .D(w25));   //: @(537, 202) /sz:(53, 64) /sn:0 /p:[ Ti0>41 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g312 (w224) @(1353, 3058) /w:[ -1 2 1 4 ]
  //: joint g262 (w198) @(739, 2631) /w:[ -1 2 1 4 ]
  //: joint g149 (w104) @(363, 1612) /w:[ 8 7 -1 10 ]
  //: joint g338 (w30) @(702, 185) /w:[ -1 2 1 4 ]
  INV1 g301 (.in(w236), .out(w260));   //: @(366, 3267) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>33 Bo0<0 ]
  assign w238 = B[6]; //: TAP g286 @(866,3025) /sn:0 /R:1 /w:[ 1 133 134 ] /ss:1
  FS g207 (.B(w174), .A(w160), .Bin(w176), .Bout(w173), .D(w178));   //: @(704, 2242) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  assign w252 = B[1]; //: TAP g296 @(1288,3025) /sn:0 /R:1 /w:[ 1 143 144 ] /ss:1
  FS g48 (.A(w34), .B(w44), .Bin(w49), .Bout(w46), .D(w51));   //: @(535, 577) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  MUX2 g200 (.in1(w164), .in0(w167), .c(w137), .out(w169));   //: @(1020, 2136) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>27 Bo0<3 ]
  MUX2 g276 (.in1(w199), .in0(w223), .c(w201), .out(w234));   //: @(1149, 2931) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>25 Bo0<3 ]
  MUX2 g29 (.in0(w13), .in1(w31), .c(w3), .out(w42));   //: @(310, 339) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>13 Li0>19 Bo0<3 ]
  //: joint g25 (w31) @(473, 174) /w:[ 7 -1 8 34 ]
  assign w16 = B[3]; //: TAP g17 @(496,127) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  //: joint g271 (w204) @(986, 2636) /w:[ -1 2 1 4 ]
  //: joint g106 (w70) @(748, 995) /w:[ -1 2 1 4 ]
  MUX2 g273 (.in1(w197), .in0(w220), .c(w201), .out(w233));   //: @(1064, 2904) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>21 Bo0<3 ]
  //: joint g83 (w97) @(144, 900) /w:[ 24 23 -1 26 ]
  assign w142 = B[5]; //: TAP g174 @(639,1804) /sn:0 /R:1 /w:[ 0 77 78 ] /ss:1
  //: GROUND g300 (w258) @(1410,3084) /sn:0 /R:2 /w:[ 0 ]
  assign w84 = B[1]; //: TAP g100 @(773,967) /sn:0 /R:1 /w:[ 0 49 50 ] /ss:1
  //: joint g193 (w134) @(785, 1830) /w:[ 2 1 4 -1 ]
  //: joint g80 (w36) @(715, 567) /w:[ -1 2 1 4 ]
  MUX2 g329 (.in1(w235), .in0(w256), .c(w236), .out(w276));   //: @(1261, 3364) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>3 Bo0<1 ]
  assign w75 = B[4]; //: TAP g94 @(512,967) /sn:0 /R:1 /w:[ 0 43 44 ] /ss:1
  //: joint g202 (w137) @(254, 2135) /w:[ 24 23 -1 26 ]
  FS g248 (.B(w207), .A(w200), .Bin(w209), .Bout(w206), .D(w211));   //: @(806, 2649) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>0 Lo0<0 Bo0<0 ]
  assign w213 = B[3]; //: TAP g253 @(1011,2605) /sn:0 /R:1 /w:[ 1 121 122 ] /ss:1
  //: joint g159 (w103) @(865, 1401) /w:[ -1 2 1 4 ]
  MUX2 g270 (.in1(w204), .in0(w217), .c(w201), .out(w232));   //: @(984, 2876) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>17 Bo0<3 ]
  //: joint g21 (w31) @(143, 174) /w:[ 19 -1 20 22 ]
  assign w125 = B[7]; //: TAP g172 @(474,1804) /sn:0 /R:1 /w:[ 0 73 74 ] /ss:1
  //: joint g232 (w170) @(246, 2399) /w:[ 2 28 -1 1 ]
  //: joint g155 (w102) @(773, 1402) /w:[ -1 2 1 4 ]
  //: joint g41 (w31) @(472, 189) /w:[ -1 35 36 38 ]
  assign w123 = A[4]; //: TAP g141 @(1360,584) /sn:0 /R:2 /w:[ 3 8 7 ] /ss:0
  FS g256 (.B(w219), .A(w199), .Bin(w221), .Bout(w218), .D(w223));   //: @(1138, 2653) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  FS g291 (.B(w246), .A(w233), .Bin(w248), .Bout(w245), .D(w250));   //: @(1075, 3075) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>0 Lo0<0 Bo0<0 ]
  FS g287 (.B(w240), .A(w231), .Bin(w242), .Bout(w239), .D(w244));   //: @(910, 3073) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g123 (B) @(1039, 1374) /w:[ -1 53 54 148 ]
  MUX2 g151 (.in0(w118), .in1(w101), .c(w104), .out(w133));   //: @(685, 1654) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>17 Bo0<3 ]
  assign w61 = B[6]; //: TAP g90 @(347,967) /sn:0 /R:1 /w:[ 0 39 40 ] /ss:1
  MUX2 g222 (.in1(w156), .in0(w175), .c(w170), .out(w196));   //: @(632, 2378) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>5 Bo0<1 ]
  MUX2 g82 (.in0(w60), .in1(w56), .c(w97), .out(w70));   //: @(798, 904) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>27 Bo0<3 ]
  FS g128 (.A(w100), .B(w108), .Bin(w113), .Bout(w110), .D(w115));   //: @(580, 1415) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g243 (B) @(283, 2206) /w:[ 92 -1 91 110 ]
  FS g91 (.A(w66), .B(w73), .Bin(w77), .Bout(w74), .D(w79));   //: @(392, 1004) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g33 (.in0(w21), .in1(w31), .c(w3), .out(w26));   //: @(482, 385) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>37 Li0>11 Bo0<3 ]
  //: joint g269 (w202) @(901, 2636) /w:[ -1 2 1 4 ]
  FS g49 (.A(w35), .B(w47), .Bin(w52), .Bout(w49), .D(w54));   //: @(619, 578) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w108 = B[4]; //: TAP g137 @(618,1372) /sn:0 /R:1 /w:[ 0 64 63 ] /ss:1
  //: joint g198 (w137) @(254, 2112) /w:[ 20 19 -1 22 ]
  FS g51 (.A(w56), .B(w53), .Bin(w59), .Bout(w55), .D(w60));   //: @(796, 580) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  //: joint g158 (w104) @(363, 1706) /w:[ 20 19 -1 22 ]
  FS g89 (.A(w65), .B(w61), .Bin(w74), .Bout(w62), .D(w76));   //: @(308, 1003) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FS g217 (.B(w189), .A(w140), .Bin(w192), .Bout(w188), .D(w193));   //: @(1116, 2247) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g77 (w35) @(632, 565) /w:[ -1 2 1 4 ]
  INV1 g302 (.in(w201), .out(w261));   //: @(311, 3267) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  FS g2 (.A(w31), .B(w0), .Bin(w2), .Bout(w3), .D(w4));   //: @(130, 197) /sz:(53, 64) /sn:0 /p:[ Ti0>23 Ti1>1 Ri0>1 Lo0<27 Bo0<1 ]
  assign w243 = B[4]; //: TAP g290 @(1033,3025) /sn:0 /R:1 /w:[ 1 137 138 ] /ss:1
  MUX2 g148 (.in0(w115), .in1(w100), .c(w104), .out(w131));   //: @(596, 1625) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>13 Bo0<3 ]
  FS g213 (.B(w183), .A(w168), .Bin(w185), .Bout(w182), .D(w187));   //: @(951, 2245) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  FS g252 (.B(w213), .A(w204), .Bin(w215), .Bout(w212), .D(w217));   //: @(973, 2651) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g72 (w97) @(144, 792) /w:[ 8 7 -1 10 ]
  FS g203 (.B(w144), .A(w152), .Bin(w148), .Bout(w170), .D(w171));   //: @(537, 2240) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<29 Bo0<0 ]
  FS g99 (.A(w70), .B(w84), .Bin(w89), .Bout(w86), .D(w91));   //: @(735, 1008) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g161 (w104) @(363, 1736) /w:[ 24 23 -1 26 ]
  MUX2 g182 (.in1(w18), .in0(w132), .c(w137), .out(w152));   //: @(527, 1985) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>5 Bo0<1 ]
  //: joint g196 (w137) @(254, 2086) /w:[ 16 15 -1 18 ]
  //: joint g189 (w133) @(709, 1831) /w:[ -1 2 4 1 ]
  //: joint g152 (w101) @(682, 1397) /w:[ -1 2 1 4 ]
  //: joint g103 (w90) @(836, 992) /w:[ -1 2 1 4 ]
  FS g246 (.B(w205), .A(w198), .Bin(w206), .Bout(w195), .D(w208));   //: @(726, 2648) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  assign w216 = B[2]; //: TAP g255 @(1091,2605) /sn:0 /R:1 /w:[ 1 123 124 ] /ss:1
  assign w240 = B[5]; //: TAP g288 @(949,3025) /sn:0 /R:1 /w:[ 1 135 136 ] /ss:1
  //: GROUND g10 (w32) @(798,208) /sn:0 /R:2 /w:[ 0 ]
  assign w180 = B[3]; //: TAP g212 @(904,2204) /sn:0 /R:1 /w:[ 1 101 102 ] /ss:1
  //: joint g199 (w136) @(942, 1834) /w:[ -1 2 1 4 ]
  assign D = {w267, w266, w265, w264, w263, w262, w261, w260}; //: CONCAT g309  @(194,3417) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g32 (w3) @(206, 362) /w:[ 18 20 -1 17 ]
  MUX2 g27 (.in0(w9), .in1(w31), .c(w3), .out(w14));   //: @(228, 316) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>17 Li0>23 Bo0<1 ]
  MUX2 g102 (.in0(w76), .in1(w65), .c(w71), .out(w95));   //: @(319, 1142) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>5 Bo0<0 ]
  //: joint g187 (w137) @(254, 2008) /w:[ 4 -1 3 6 ]
  MUX2 g240 (.in1(w140), .in0(w193), .c(w170), .out(w199));   //: @(1127, 2552) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>27 Bo0<3 ]
  assign w39 = B[5]; //: TAP g57 @(407,542) /sn:0 /R:1 /w:[ 0 30 29 ] /ss:1
  FS g9 (.A(w30), .B(w28), .Bin(w32), .Bout(w27), .D(w33));   //: @(689, 204) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g71 (w26) @(462, 563) /w:[ -1 2 1 4 ]
  MUX2 g142 (.in0(w109), .in1(w98), .c(w104), .out(w130));   //: @(421, 1560) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>5 Bo0<0 ]
  //: joint g318 (w236) @(633, 3258) /w:[ 22 24 -1 21 ]
  assign w255 = B[0]; //: TAP g298 @(1379,3025) /sn:0 /R:1 /w:[ 1 145 146 ] /ss:1
  FS g295 (.B(w252), .A(w235), .Bin(w254), .Bout(w251), .D(w256));   //: @(1250, 3077) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g145 (w99) @(504, 1397) /w:[ -1 2 1 4 ]
  //: joint g327 (w236) @(633, 3343) /w:[ 10 12 -1 9 ]
  MUX2 g73 (.in0(w51), .in1(w34), .c(w97), .out(w96));   //: @(551, 823) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>17 Bo0<3 ]
  //: GROUND g180 (w128) @(1084,1859) /sn:0 /R:2 /w:[ 0 ]
  //: joint g42 (w3) @(206, 456) /w:[ 2 4 -1 1 ]
  //: joint g74 (w34) @(548, 563) /w:[ -1 2 1 4 ]
  assign w224 = A[0]; //: TAP g299 @(1360,2820) /sn:0 /R:2 /w:[ 3 16 15 ] /ss:0
  assign w164 = A[3]; //: TAP g181 @(1360,740) /sn:0 /R:2 /w:[ 3 10 9 ] /ss:0
  FS g168 (.A(w134), .B(w150), .Bin(w153), .Bout(w149), .D(w155));   //: @(762, 1848) /sz:(53, 64) /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  MUX2 g79 (.in0(w57), .in1(w36), .c(w97), .out(w69));   //: @(724, 877) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>25 Bo0<3 ]
  MUX2 g117 (.in0(w91), .in1(w70), .c(w71), .out(w102));   //: @(753, 1271) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>25 Bo0<3 ]
  MUX2 g194 (.in1(w135), .in0(w159), .c(w137), .out(w166));   //: @(855, 2089) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>21 Bo0<3 ]
  FS g215 (.B(w186), .A(w169), .Bin(w188), .Bout(w185), .D(w190));   //: @(1031, 2246) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g36 (w3) @(206, 408) /w:[ 10 12 -1 9 ]
  assign w186 = B[1]; //: TAP g216 @(1069,2204) /sn:0 /R:1 /w:[ 1 105 106 ] /ss:1
  assign w158 = B[1]; //: TAP g178 @(968,1804) /sn:0 /R:1 /w:[ 0 85 86 ] /ss:1
  MUX2 g144 (.in0(w112), .in1(w99), .c(w104), .out(w18));   //: @(508, 1589) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>9 Bo0<3 ]
  assign w64 = B[7]; //: TAP g125 @(367,1372) /sn:0 /R:1 /w:[ 0 70 69 ] /ss:1
  //: joint g81 (w97) @(144, 874) /w:[ 20 19 -1 22 ]
  //: joint g275 (w197) @(1066, 2630) /w:[ -1 2 1 4 ]
  //: joint g22 (w31) @(230, 174) /w:[ 15 16 18 24 ]
  FS g45 (.A(w42), .B(w6), .Bin(w40), .Bout(w10), .D(w257));   //: @(287, 574) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  MUX2 g70 (.in0(w48), .in1(w26), .c(w97), .out(w66));   //: @(466, 797) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>13 Bo0<3 ]
  //: joint g282 (B) @(302, 2607) /w:[ 112 -1 111 130 ]
  MUX2 g114 (.in0(w88), .in1(w69), .c(w71), .out(w101));   //: @(661, 1248) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Li0>21 Bo0<3 ]
  FS g209 (.B(w177), .A(w165), .Bin(w179), .Bout(w176), .D(w181));   //: @(784, 2243) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g229 (w166) @(879, 2226) /w:[ -1 2 1 4 ]
  MUX2 g279 (.in1(w191), .in0(w226), .c(w201), .out(w235));   //: @(1239, 2963) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>27 Bo0<3 ]
  MUX2 g323 (.in1(w233), .in0(w250), .c(w236), .out(w274));   //: @(1086, 3320) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Li0>11 Bo0<1 ]
  FS g164 (.A(w130), .B(w125), .Bin(w129), .Bout(w137), .D(w138));   //: @(434, 1844) /sz:(53, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<29 Bo0<1 ]
  //: joint g30 (w3) @(206, 333) /w:[ 22 -1 24 21 ]
  //: joint g118 (w66) @(405, 990) /w:[ -1 2 1 4 ]
  FS g289 (.B(w243), .A(w232), .Bin(w245), .Bout(w242), .D(w247));   //: @(995, 3074) /sz:(53, 64) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>1 Lo0<0 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin HA
module HA(Cout, S, B, A);
//: interface  /sz:(40, 54) /bd:[ Ti0>B(29/40) Ti1>A(10/40) Lo0<Cout(32/54) Bo0<S(21/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(180,139)(165,139)(165,230){1}
//: {2}(167,232)(198,232){3}
//: {4}(163,232)(92,232){5}
input A;    //: /sn:0 {0}(198,212)(142,212)(142,123){1}
//: {2}(144,121)(180,121){3}
//: {4}(140,121)(97,121){5}
output Cout;    //: /sn:0 {0}(329,221)(255,221)(255,221)(240,221){1}
output S;    //: /sn:0 {0}(328,138)(253,138)(253,138)(237,138){1}
//: enddecls

  EXOR2 g4 (.a(A), .b(B), .out(S));   //: @(181, 111) /sz:(55, 42) /sn:0 /p:[ Li0>3 Li1>0 Ro0<1 ]
  //: OUT g3 (Cout) @(326,221) /sn:0 /w:[ 0 ]
  //: OUT g2 (S) @(325,138) /sn:0 /w:[ 0 ]
  //: IN g1 (B) @(90,232) /sn:0 /w:[ 5 ]
  //: joint g6 (B) @(165, 232) /w:[ 2 1 4 -1 ]
  //: joint g7 (A) @(142, 121) /w:[ 2 -1 4 1 ]
  AND2 g5 (.in1(A), .in2(B), .out(Cout));   //: @(199, 202) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>3 Ro0<1 ]
  //: IN g0 (A) @(95,121) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin REG8sINaddsub
module REG8sINaddsub(mode, ctrl, out, Out2, clk, in);
//: interface  /sz:(56, 117) /bd:[ Ti0>in[7:0](24/56) Li0>clk(78/117) Li1>ctrl(39/117) Ri0>mode(39/117) Bo0<out(24/56) Ro0<Out2[7:0](97/117) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] in;    //: /sn:0 {0}(#:21,25)(21,33)(22,33)(22,47){1}
//: {2}(22,48)(22,183){3}
//: {4}(22,184)(22,317){5}
//: {6}(22,318)(22,453){7}
//: {8}(22,454)(22,601){9}
//: {10}(22,602)(22,740){11}
//: {12}(22,741)(22,868){13}
//: {14}(22,869)(22,1030){15}
//: {16}(22,1031)(22,1048){17}
output out;    //: /sn:0 {0}(508,1049)(531,1049){1}
//: {2}(535,1049)(552,1049){3}
//: {4}(533,1047)(533,1025)(786,1025)(786,485)(978,485){5}
supply0 w3;    //: /sn:0 {0}(301,43)(322,43)(322,36)(343,36){1}
output [7:0] Out2;    //: /sn:0 {0}(1037,450)(#:984,450){1}
input mode;    //: /sn:0 {0}(222,71)(222,125)(604,125)(604,289){1}
//: {2}(602,291)(225,291)(225,211){3}
//: {4}(604,293)(604,428){5}
//: {6}(602,430)(224,430)(224,344){7}
//: {8}(604,432)(604,572){9}
//: {10}(602,574)(227,574)(227,481){11}
//: {12}(604,576)(604,710){13}
//: {14}(602,712)(228,712)(228,629){15}
//: {16}(604,714)(604,834){17}
//: {18}(602,836)(233,836)(233,768){19}
//: {20}(604,838)(604,991){21}
//: {22}(602,993)(234,993)(234,898){23}
//: {24}(604,995)(604,1141){25}
//: {26}(602,1143)(236,1143)(236,1059){27}
//: {28}(604,1145)(604,1157){29}
input ctrl;    //: /sn:0 {0}(363,206)(363,285)(639,285){1}
//: {2}(641,283)(641,118)(361,118)(361,70){3}
//: {4}(641,287)(641,422){5}
//: {6}(639,424)(365,424)(365,342){7}
//: {8}(641,426)(641,567){9}
//: {10}(639,569)(365,569)(365,484){11}
//: {12}(641,571)(641,704){13}
//: {14}(639,706)(365,706)(365,627){15}
//: {16}(641,708)(641,829){17}
//: {18}(639,831)(366,831)(366,766){19}
//: {20}(641,833)(641,985){21}
//: {22}(639,987)(365,987)(365,898){23}
//: {24}(641,989)(641,1134){25}
//: {26}(639,1136)(364,1136)(364,1060){27}
//: {28}(641,1138)(641,1157){29}
input clk;    //: /sn:0 {0}(482,217)(482,278)(677,278){1}
//: {2}(679,276)(679,140)(486,140)(486,81){3}
//: {4}(679,280)(679,411){5}
//: {6}(677,413)(482,413)(482,353){7}
//: {8}(679,415)(679,557){9}
//: {10}(677,559)(483,559)(483,495){11}
//: {12}(679,561)(679,695){13}
//: {14}(677,697)(486,697)(486,638){15}
//: {16}(679,699)(679,818){17}
//: {18}(677,820)(485,820)(485,777){19}
//: {20}(679,822)(679,976){21}
//: {22}(677,978)(484,978)(484,909){23}
//: {24}(679,980)(679,1122){25}
//: {26}(677,1124)(485,1124)(485,1071){27}
//: {28}(679,1126)(679,1158){29}
wire w6;    //: /sn:0 {0}(135,76)(169,76)(169,56)(204,56){1}
wire w32;    //: /sn:0 {0}(347,308)(337,308)(337,289)(531,289)(531,223){1}
//: {2}(533,221)(957,221)(957,425)(978,425){3}
//: {4}(531,219)(531,195)(505,195){5}
wire w7;    //: /sn:0 {0}(467,59)(412,59)(412,45)(385,45){1}
wire w60;    //: /sn:0 {0}(466,1049)(413,1049)(413,1035)(388,1035){1}
wire w16;    //: /sn:0 {0}(145,1063)(187,1063)(187,1044)(218,1044){1}
wire w15;    //: /sn:0 {0}(148,772)(186,772)(186,753)(215,753){1}
wire w4;    //: /sn:0 {0}(138,349)(172,349)(172,329)(206,329){1}
wire w0;    //: /sn:0 {0}(26,48)(72,48){1}
//: {2}(76,48)(193,48)(193,37)(204,37){3}
//: {4}(74,50)(74,77)(93,77){5}
wire w21;    //: /sn:0 {0}(348,732)(334,732)(334,709)(532,709)(532,649){1}
//: {2}(534,647)(719,647)(719,455)(978,455){3}
//: {4}(532,645)(532,616)(509,616){5}
wire w58;    //: /sn:0 {0}(260,1034)(303,1034)(303,1045)(346,1045){1}
wire w31;    //: /sn:0 {0}(347,450)(335,450)(335,429)(532,429)(532,370){1}
//: {2}(534,368)(949,368)(949,435)(978,435){3}
//: {4}(532,366)(532,331)(505,331){5}
wire w28;    //: /sn:0 {0}(464,473)(412,473)(412,459)(389,459){1}
wire w41;    //: /sn:0 {0}(26,741)(75,741){1}
//: {2}(79,741)(147,741)(147,734)(215,734){3}
//: {4}(77,743)(77,773)(106,773){5}
wire w23;    //: /sn:0 {0}(26,602)(72,602){1}
//: {2}(76,602)(143,602)(143,595)(210,595){3}
//: {4}(74,604)(74,634)(105,634){5}
wire w36;    //: /sn:0 {0}(467,616)(414,616)(414,602)(389,602){1}
wire w20;    //: /sn:0 {0}(463,331)(412,331)(412,317)(389,317){1}
wire w24;    //: /sn:0 {0}(347,864)(332,864)(332,834)(533,834)(533,793){1}
//: {2}(535,791)(734,791)(734,465)(978,465){3}
//: {4}(533,789)(533,755)(508,755){5}
wire w1;    //: /sn:0 {0}(139,216)(173,216)(173,196)(207,196){1}
wire w25;    //: /sn:0 {0}(252,604)(304,604)(304,612)(347,612){1}
wire w18;    //: /sn:0 {0}(248,319)(304,319)(304,327)(347,327){1}
wire w8;    //: /sn:0 {0}(249,186)(302,186)(302,191)(345,191){1}
wire w30;    //: /sn:0 {0}(978,445)(704,445)(704,504)(533,504){1}
//: {2}(531,502)(531,473)(506,473){3}
//: {4}(531,506)(531,573)(332,573)(332,593)(347,593){5}
wire w12;    //: /sn:0 {0}(156,903)(186,903)(186,883)(216,883){1}
wire w11;    //: /sn:0 {0}(147,633)(176,633)(176,614)(210,614){1}
wire w57;    //: /sn:0 {0}(26,1031)(79,1031){1}
//: {2}(83,1031)(156,1031)(156,1025)(218,1025){3}
//: {4}(81,1033)(81,1064)(103,1064){5}
wire w49;    //: /sn:0 {0}(26,869)(76,869){1}
//: {2}(80,869)(154,869)(154,864)(216,864){3}
//: {4}(78,871)(78,904)(114,904){5}
wire w44;    //: /sn:0 {0}(466,755)(414,755)(414,741)(390,741){1}
wire w2;    //: /sn:0 {0}(26,184)(74,184){1}
//: {2}(78,184)(142,184)(142,177)(207,177){3}
//: {4}(76,186)(76,217)(97,217){5}
wire w10;    //: /sn:0 {0}(463,195)(411,195)(411,181)(387,181){1}
wire w13;    //: /sn:0 {0}(26,318)(76,318){1}
//: {2}(80,318)(198,318)(198,310)(206,310){3}
//: {4}(78,320)(78,350)(96,350){5}
wire w27;    //: /sn:0 {0}(346,1026)(335,1026)(335,993)(534,993)(534,927){1}
//: {2}(536,925)(753,925)(753,475)(978,475){3}
//: {4}(534,923)(534,887)(507,887){5}
wire w52;    //: /sn:0 {0}(465,887)(413,887)(413,873)(389,873){1}
wire w5;    //: /sn:0 {0}(246,46)(300,46)(300,55)(343,55){1}
wire w33;    //: /sn:0 {0}(345,172)(335,172)(335,152)(519,152)(519,95){1}
//: {2}(521,93)(963,93)(963,415)(978,415){3}
//: {4}(519,91)(519,59)(509,59){5}
wire w29;    //: /sn:0 {0}(26,454)(71,454){1}
//: {2}(75,454)(142,454)(142,447)(209,447){3}
//: {4}(73,456)(73,488)(94,488){5}
wire w9;    //: /sn:0 {0}(136,487)(181,487)(181,466)(209,466){1}
wire w50;    //: /sn:0 {0}(258,873)(304,873)(304,883)(347,883){1}
wire w42;    //: /sn:0 {0}(257,743)(305,743)(305,751)(348,751){1}
wire w26;    //: /sn:0 {0}(251,456)(299,456)(299,469)(347,469){1}
//: enddecls

  //: joint g4 (w0) @(74, 48) /w:[ 2 -1 1 4 ]
  //: joint g61 (ctrl) @(641, 987) /w:[ -1 21 22 24 ]
  MUX2 g8 (.in0(w2), .in1(w1), .c(mode), .out(w8));   //: @(208, 168) /sz:(40, 42) /sn:0 /p:[ Li0>3 Li1>1 Bi0>3 Ro0<0 ]
  //: joint g37 (w41) @(77, 741) /w:[ 2 -1 1 4 ]
  //: joint g58 (mode) @(604, 291) /w:[ -1 1 2 4 ]
  //: joint g55 (mode) @(604, 712) /w:[ -1 13 14 16 ]
  //: IN g51 (mode) @(604,1159) /sn:0 /R:1 /w:[ 29 ]
  MUX2 g34 (.in0(w41), .in1(w15), .c(mode), .out(w42));   //: @(216, 725) /sz:(40, 42) /sn:0 /p:[ Li0>3 Li1>1 Bi0>19 Ro0<0 ]
  FFD g13 (.D(w10), .Clk(clk), .Y(w32));   //: @(464, 176) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>0 Ro0<5 ]
  assign w0 = in[7]; //: TAP g3 @(20,48) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: joint g65 (ctrl) @(641, 424) /w:[ -1 5 6 8 ]
  MUX2 g2 (.in0(w0), .in1(w6), .c(mode), .out(w5));   //: @(205, 28) /sz:(40, 42) /sn:0 /p:[ Li0>3 Li1>1 Bi0>0 Ro0<0 ]
  assign Out2 = {w33, w32, w31, w30, w21, w24, w27, out}; //: CONCAT g76  @(983,450) /sn:0 /w:[ 1 3 3 3 0 3 3 3 5 ] /dr:0 /tp:0 /drp:1
  //: joint g77 (w33) @(519, 93) /w:[ 2 4 -1 1 ]
  //: IN g59 (ctrl) @(641,1159) /sn:0 /R:1 /w:[ 29 ]
  //: joint g72 (clk) @(679, 559) /w:[ -1 9 10 12 ]
  INV1 g1 (.in(w0), .out(w6));   //: @(94, 56) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g64 (ctrl) @(641, 569) /w:[ -1 9 10 12 ]
  //: joint g11 (w2) @(76, 184) /w:[ 2 -1 1 4 ]
  MUX2 g16 (.in0(w13), .in1(w4), .c(mode), .out(w18));   //: @(207, 301) /sz:(40, 42) /sn:0 /p:[ Li0>3 Li1>1 Bi0>7 Ro0<0 ]
  //: OUT g50 (out) @(549,1049) /sn:0 /w:[ 3 ]
  MUX2 g28 (.in0(w23), .in1(w11), .c(mode), .out(w25));   //: @(211, 586) /sz:(40, 42) /sn:0 /p:[ Li0>3 Li1>1 Bi0>15 Ro0<0 ]
  assign w2 = in[6]; //: TAP g10 @(20,184) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g78 (w32) @(531, 221) /w:[ 2 4 -1 1 ]
  //: joint g19 (w13) @(78, 318) /w:[ 2 -1 1 4 ]
  MUX2 g32 (.in0(w21), .in1(w42), .c(ctrl), .out(w44));   //: @(349, 723) /sz:(40, 42) /sn:0 /p:[ Li0>0 Li1>1 Bi0>19 Ro0<1 ]
  FFD g27 (.D(w36), .Clk(clk), .Y(w21));   //: @(468, 597) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>15 Ro0<5 ]
  //: joint g69 (clk) @(679, 978) /w:[ -1 21 22 24 ]
  MUX2 g38 (.in0(w24), .in1(w50), .c(ctrl), .out(w52));   //: @(348, 855) /sz:(40, 42) /sn:0 /p:[ Li0>0 Li1>1 Bi0>23 Ro0<1 ]
  //: GROUND g6 (w3) @(295,43) /sn:0 /R:3 /w:[ 0 ]
  //: joint g57 (mode) @(604, 430) /w:[ -1 5 6 8 ]
  //: joint g53 (mode) @(604, 993) /w:[ -1 21 22 24 ]
  INV1 g9 (.in(w2), .out(w1));   //: @(98, 196) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  MUX2 g7 (.in0(w33), .in1(w8), .c(ctrl), .out(w10));   //: @(346, 163) /sz:(40, 42) /sn:0 /p:[ Li0>0 Li1>1 Bi0>0 Ro0<1 ]
  //: OUT g75 (Out2) @(1034,450) /sn:0 /w:[ 0 ]
  //: joint g31 (w23) @(74, 602) /w:[ 2 -1 1 4 ]
  //: joint g71 (clk) @(679, 697) /w:[ -1 13 14 16 ]
  MUX2 g20 (.in0(w31), .in1(w26), .c(ctrl), .out(w28));   //: @(348, 441) /sz:(40, 42) /sn:0 /p:[ Li0>0 Li1>1 Bi0>11 Ro0<1 ]
  FFD g15 (.D(w20), .Clk(clk), .Y(w31));   //: @(464, 312) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>7 Ro0<5 ]
  //: joint g68 (clk) @(679, 1124) /w:[ -1 25 26 28 ]
  //: IN g67 (clk) @(679,1160) /sn:0 /R:1 /w:[ 29 ]
  FFD g39 (.D(w52), .Clk(clk), .Y(w27));   //: @(466, 868) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>23 Ro0<5 ]
  //: joint g43 (w49) @(78, 869) /w:[ 2 -1 1 4 ]
  assign w57 = in[0]; //: TAP g48 @(20,1031) /sn:0 /R:2 /w:[ 0 16 15 ] /ss:1
  //: joint g25 (w29) @(73, 454) /w:[ 2 -1 1 4 ]
  //: joint g73 (clk) @(679, 413) /w:[ -1 5 6 8 ]
  //: joint g62 (ctrl) @(641, 831) /w:[ -1 17 18 20 ]
  INV1 g29 (.in(w23), .out(w11));   //: @(106, 613) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  INV1 g17 (.in(w13), .out(w4));   //: @(97, 329) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g63 (ctrl) @(641, 706) /w:[ -1 13 14 16 ]
  //: joint g52 (mode) @(604, 1143) /w:[ -1 25 26 28 ]
  assign w49 = in[1]; //: TAP g42 @(20,869) /sn:0 /R:2 /w:[ 0 14 13 ] /ss:1
  //: joint g83 (w27) @(534, 925) /w:[ 2 4 -1 1 ]
  //: joint g74 (clk) @(679, 278) /w:[ -1 2 1 4 ]
  //: joint g56 (mode) @(604, 574) /w:[ -1 9 10 12 ]
  MUX2 g14 (.in0(w32), .in1(w18), .c(ctrl), .out(w20));   //: @(348, 299) /sz:(40, 42) /sn:0 /p:[ Li0>0 Li1>1 Bi0>7 Ro0<1 ]
  MUX2 g5 (.in0(w3), .in1(w5), .c(ctrl), .out(w7));   //: @(344, 27) /sz:(40, 42) /sn:0 /p:[ Li0>1 Li1>1 Bi0>3 Ro0<1 ]
  INV1 g47 (.in(w57), .out(w16));   //: @(104, 1043) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  MUX2 g44 (.in0(w27), .in1(w58), .c(ctrl), .out(w60));   //: @(347, 1017) /sz:(40, 42) /sn:0 /p:[ Li0>0 Li1>1 Bi0>27 Ro0<1 ]
  //: joint g79 (w31) @(532, 368) /w:[ 2 4 -1 1 ]
  //: joint g80 (w30) @(531, 504) /w:[ 1 2 -1 4 ]
  assign w41 = in[2]; //: TAP g36 @(20,741) /sn:0 /R:2 /w:[ 0 12 11 ] /ss:1
  assign w29 = in[4]; //: TAP g24 @(20,454) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  FFD g21 (.D(w28), .Clk(clk), .Y(w30));   //: @(465, 454) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>11 Ro0<3 ]
  //: joint g84 (out) @(533, 1049) /w:[ 2 4 1 -1 ]
  INV1 g41 (.in(w49), .out(w12));   //: @(115, 883) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  INV1 g23 (.in(w29), .out(w9));   //: @(95, 467) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g60 (ctrl) @(641, 1136) /w:[ -1 25 26 28 ]
  //: joint g54 (mode) @(604, 836) /w:[ -1 17 18 20 ]
  MUX2 g40 (.in0(w49), .in1(w12), .c(mode), .out(w50));   //: @(217, 855) /sz:(40, 42) /sn:0 /p:[ Li0>3 Li1>1 Bi0>23 Ro0<0 ]
  //: joint g81 (w21) @(532, 647) /w:[ 2 4 -1 1 ]
  //: joint g70 (clk) @(679, 820) /w:[ -1 17 18 20 ]
  MUX2 g46 (.in0(w57), .in1(w16), .c(mode), .out(w58));   //: @(219, 1016) /sz:(40, 42) /sn:0 /p:[ Li0>3 Li1>1 Bi0>27 Ro0<0 ]
  FFD g45 (.D(w60), .Clk(clk), .Y(out));   //: @(467, 1030) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>27 Ro0<0 ]
  INV1 g35 (.in(w41), .out(w15));   //: @(107, 752) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  MUX2 g26 (.in0(w30), .in1(w25), .c(ctrl), .out(w36));   //: @(348, 584) /sz:(40, 42) /sn:0 /p:[ Li0>5 Li1>1 Bi0>15 Ro0<1 ]
  MUX2 g22 (.in0(w29), .in1(w9), .c(mode), .out(w26));   //: @(210, 438) /sz:(40, 42) /sn:0 /p:[ Li0>3 Li1>1 Bi0>11 Ro0<0 ]
  //: IN g0 (in) @(21,23) /sn:0 /R:3 /w:[ 0 ]
  //: joint g66 (ctrl) @(641, 285) /w:[ -1 2 1 4 ]
  //: joint g82 (w24) @(533, 791) /w:[ 2 4 -1 1 ]
  assign w13 = in[5]; //: TAP g18 @(20,318) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  FFD g12 (.D(w7), .Clk(clk), .Y(w33));   //: @(468, 40) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>3 Ro0<5 ]
  FFD g33 (.D(w44), .Clk(clk), .Y(w24));   //: @(467, 736) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>19 Ro0<5 ]
  assign w23 = in[3]; //: TAP g30 @(20,602) /sn:0 /R:2 /w:[ 0 10 9 ] /ss:1
  //: joint g49 (w57) @(81, 1031) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin Calcolatrice_4_operazioni
module Calcolatrice_4_operazioni(AxB, A, RestoDiv, Neg, Carica, Clk, AddSub, B, AdivB);
//: interface  /sz:(200, 109) /bd:[ Ti0>B[7:0](152/200) Ti1>A[7:0](40/200) Li0>Clk(22/109) Li1>Neg(71/109) Ri0>Carica(25/109) Bo0<AxB[15:0](106/200) Bo1<AddSub[8:0](42/200) Bo2<AdivB[7:0](171/200) Ro0<RestoDiv[7:0](81/109) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:243,127)(243,163){1}
output [7:0] RestoDiv;    //: /sn:0 {0}(#:582,361)(582,332)(#:613,332){1}
output [8:0] AddSub;    //: /sn:0 {0}(#:226,285)(226,245){1}
input [7:0] A;    //: /sn:0 {0}(#:164,148)(201,148)(201,163){1}
output [7:0] AdivB;    //: /sn:0 {0}(#:557,307)(557,292)(#:613,292){1}
output [15:0] AxB;    //: /sn:0 {0}(422,341)(422,310)(#:459,310){1}
input Clk;    //: /sn:0 {0}(125,227)(188,227){1}
input Neg;    //: /sn:0 {0}(376,59)(376,46)(439,46){1}
//: {2}(441,44)(441,34){3}
//: {4}(441,48)(441,186)(263,186){5}
input Carica;    //: /sn:0 {0}(357,127)(357,70)(110,70){1}
//: {2}(106,70)(90,70)(90,187)(64,187){3}
//: {4}(108,72)(108,185)(188,185){5}
wire [7:0] w6;    //: /sn:0 {0}(#:263,214)(320,214)(320,201)(#:335,201){1}
wire [7:0] w0;    //: /sn:0 {0}(#:400,201)(507,201)(507,212){1}
//: {2}(509,214)(662,214)(#:662,271){3}
//: {4}(507,216)(507,228)(508,228)(#:508,277){5}
wire [7:0] w3;    //: /sn:0 {0}(#:400,249)(468,249)(468,250)(478,250){1}
//: {2}(480,248)(480,236)(632,236)(#:632,271){3}
//: {4}(480,252)(#:480,277){5}
wire w1;    //: /sn:0 {0}(368,169)(368,184){1}
wire [7:0] w2;    //: /sn:0 {0}(#:263,238)(320,238)(320,249)(#:335,249){1}
wire w5;    //: /sn:0 {0}(377,101)(377,118)(377,118)(377,127){1}
//: enddecls

  //: OUT g8 (AxB) @(422,338) /sn:0 /R:3 /w:[ 0 ]
  //: IN g4 (A) @(162,148) /sn:0 /w:[ 0 ]
  //: OUT g13 (RestoDiv) @(582,358) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (Neg) @(441,32) /sn:0 /R:3 /w:[ 3 ]
  //: IN g2 (Carica) @(62,187) /sn:0 /w:[ 3 ]
  //: IN g1 (Clk) @(123,227) /sn:0 /w:[ 0 ]
  INV1 g16 (.in(Neg), .out(w5));   //: @(357, 60) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  AND2 g11 (.in1(w5), .in2(Carica), .out(w1));   //: @(347, 128) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<0 ]
  Mux8 g10 (.ctrl(w1), .B(w2), .A(w6), .B2(w3), .A1(w0));   //: @(336, 185) /sz:(63, 80) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: OUT g6 (AddSub) @(226,282) /sn:0 /R:3 /w:[ 0 ]
  Mul16b g7 (.B(w3), .A(w0), .S(AxB));   //: @(460, 278) /sz:(64, 63) /R:3 /sn:0 /p:[ Ti0>5 Ti1>5 Lo0<1 ]
  Div8b g9 (.B(w3), .A(w0), .R(RestoDiv), .D(AdivB));   //: @(614, 272) /sz:(64, 80) /R:3 /sn:0 /p:[ Ti0>3 Ti1>3 Lo0<1 Lo1<1 ]
  //: joint g15 (w0) @(507, 214) /w:[ 2 1 -1 4 ]
  //: joint g17 (Carica) @(108, 70) /w:[ 1 -1 2 4 ]
  //: joint g14 (w3) @(480, 250) /w:[ -1 2 1 4 ]
  //: IN g5 (B) @(243,125) /sn:0 /R:3 /w:[ 0 ]
  BySaddsub2 g0 (.B(B), .A(A), .clk(Clk), .load(Carica), .mode(Neg), .S(AddSub), .A2(w6), .B2(w2));   //: @(189, 164) /sz:(73, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Li1>5 Ri0>5 Bo0<1 Ro0<0 Ro1<0 ]
  //: joint g18 (Neg) @(441, 46) /w:[ -1 2 1 4 ]
  //: OUT g12 (AdivB) @(557,304) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin AND2
module AND2(in2, in1, out);
//: interface  /sz:(40, 40) /bd:[ Li0>in2(30/40) Li1>in1(10/40) Ro0<out(19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output out;    //: /sn:0 {0}(402,172)(415,172)(415,172)(436,172){1}
input in1;    //: /sn:0 {0}(284,165)(273,165)(273,165)(249,165){1}
input in2;    //: /sn:0 {0}(284,185)(273,185)(273,185)(249,185){1}
wire w2;    //: /sn:0 {0}(326,173)(338,173)(338,173)(360,173){1}
//: enddecls

  //: IN g4 (in2) @(247,185) /sn:0 /w:[ 1 ]
  //: IN g3 (in1) @(247,165) /sn:0 /w:[ 1 ]
  //: OUT g2 (out) @(433,172) /sn:0 /w:[ 1 ]
  INV1 g1 (.in(w2), .out(out));   //: @(361, 152) /sz:(40, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  NAND2 g0 (.in1(in1), .in2(in2), .out(w2));   //: @(285, 155) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin EXOR2
module EXOR2(out, b, a);
//: interface  /sz:(55, 42) /bd:[ Li0>b(28/42) Li1>a(10/42) Ro0<out(27/42) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(149,200)(109,200)(109,185){1}
//: {2}(111,183)(114,183)(114,167)(218,167)(218,101)(270,101){3}
//: {4}(107,183)(96,183)(96,183)(86,183){5}
output out;    //: /sn:0 {0}(439,157)(474,157)(474,157)(489,157){1}
input a;    //: /sn:0 {0}(153,82)(118,82)(118,82)(108,82){1}
//: {2}(104,82)(97,82)(97,82)(91,82){3}
//: {4}(106,84)(106,122)(227,122)(227,179)(263,179){5}
wire w6;    //: /sn:0 {0}(312,89)(382,89)(382,149)(397,149){1}
wire w3;    //: /sn:0 {0}(191,199)(248,199)(248,199)(263,199){1}
wire w1;    //: /sn:0 {0}(195,81)(255,81)(255,81)(270,81){1}
wire w9;    //: /sn:0 {0}(305,187)(382,187)(382,169)(397,169){1}
//: enddecls

  //: joint g8 (a) @(106, 82) /w:[ 1 -1 2 4 ]
  INV1 g4 (.in(b), .out(w3));   //: @(150, 179) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  INV1 g3 (.in(a), .out(w1));   //: @(154, 61) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: OUT g2 (out) @(486,157) /sn:0 /w:[ 1 ]
  //: IN g1 (b) @(84,183) /sn:0 /w:[ 5 ]
  NAND2 g6 (.in2(w3), .in1(a), .out(w9));   //: @(264, 169) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>5 Ro0<0 ]
  //: joint g9 (b) @(109, 183) /w:[ 2 -1 4 1 ]
  NAND2 g7 (.in2(w9), .in1(w6), .out(out));   //: @(398, 139) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  NAND2 g5 (.in2(b), .in1(w1), .out(w6));   //: @(271, 71) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]
  //: IN g0 (a) @(89,82) /sn:0 /w:[ 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin REG8sIN
module REG8sIN(out, in, clk, putM, ctrl);
//: interface  /sz:(49, 82) /bd:[ Ti0>clk(24/49) Li0>in[7:0](49/82) Bi0>ctrl(9/49) Bo0<out(41/49) Ro0<putM[7:0](48/82) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] in;    //: /sn:0 {0}(#:13,631)(13,622){1}
//: {2}(13,621)(13,533){3}
//: {4}(13,532)(13,437){5}
//: {6}(13,436)(13,362){7}
//: {8}(13,361)(13,289){9}
//: {10}(13,288)(13,211){11}
//: {12}(13,210)(13,126){13}
//: {14}(13,125)(13,44){15}
//: {16}(13,43)(#:13,17){17}
output out;    //: /sn:0 {0}(291,640)(250,640)(250,620){1}
//: {2}(252,618)(500,618)(500,408)(517,408){3}
//: {4}(250,616)(250,615)(235,615){5}
supply0 w25;    //: /sn:0 {0}(50,32)(80,32){1}
input ctrl;    //: /sn:0 {0}(94,637)(94,656)(373,656){1}
//: {2}(375,654)(375,551){3}
//: {4}(375,547)(375,484){5}
//: {6}(375,480)(375,391){7}
//: {8}(375,387)(375,322){9}
//: {10}(375,318)(375,238){11}
//: {12}(375,234)(375,153){13}
//: {14}(375,149)(375,85)(98,85)(98,66){15}
//: {16}(373,151)(98,151)(98,144){17}
//: {18}(373,236)(97,236)(97,227){19}
//: {20}(373,320)(93,320)(93,302){21}
//: {22}(373,389)(94,389)(94,379){23}
//: {24}(373,482)(93,482)(93,453){25}
//: {26}(373,549)(351,549)(351,582)(95,582)(95,549){27}
//: {28}(375,658)(375,683){29}
output [7:0] putM;    //: /sn:0 {0}(602,380)(538,380)(#:538,373)(#:523,373){1}
input clk;    //: /sn:0 {0}(212,637)(212,667)(324,667){1}
//: {2}(326,665)(326,562){3}
//: {4}(326,558)(326,471){5}
//: {6}(326,467)(326,397){7}
//: {8}(326,393)(326,316){9}
//: {10}(326,312)(326,244){11}
//: {12}(326,240)(326,163){13}
//: {14}(326,159)(326,78)(212,78)(212,63){15}
//: {16}(324,161)(212,161)(212,144){17}
//: {18}(324,242)(210,242)(210,225){19}
//: {20}(324,314)(211,314)(211,298){21}
//: {22}(324,395)(213,395)(213,375){23}
//: {24}(324,469)(216,469)(216,451){25}
//: {26}(324,560)(209,560)(209,545){27}
//: {28}(326,669)(326,687){29}
wire w32;    //: /sn:0 {0}(76,364)(46,364)(46,362)(17,362){1}
wire w6;    //: /sn:0 {0}(121,202)(148,202)(148,203)(191,203){1}
wire w7;    //: /sn:0 {0}(122,119)(157,119)(157,122)(193,122){1}
wire w16;    //: /sn:0 {0}(76,622)(17,622){1}
wire w14;    //: /sn:0 {0}(517,378)(456,378)(456,353)(248,353){1}
//: {2}(244,353)(236,353){3}
//: {4}(246,355)(246,404)(60,404)(60,419)(75,419){5}
wire w4;    //: /sn:0 {0}(193,615)(133,615)(133,612)(118,612){1}
wire w15;    //: /sn:0 {0}(117,428)(143,428)(143,429)(197,429){1}
wire w0;    //: /sn:0 {0}(122,41)(193,41){1}
wire w34;    //: /sn:0 {0}(75,438)(25,438)(25,437)(17,437){1}
wire w28;    //: /sn:0 {0}(79,212)(48,212)(48,211)(17,211){1}
wire w36;    //: /sn:0 {0}(77,534)(25,534)(25,533)(17,533){1}
wire w23;    //: /sn:0 {0}(80,51)(25,51)(25,44)(17,44){1}
wire w1;    //: /sn:0 {0}(76,603)(61,603)(61,573)(242,573)(242,525){1}
//: {2}(242,521)(242,513)(489,513)(489,398)(517,398){3}
//: {4}(240,523)(232,523){5}
wire w18;    //: /sn:0 {0}(119,524)(140,524)(140,523)(190,523){1}
wire w8;    //: /sn:0 {0}(517,358)(481,358)(481,203)(245,203){1}
//: {2}(241,203)(233,203){3}
//: {4}(243,205)(243,253)(60,253)(60,268)(75,268){5}
wire w30;    //: /sn:0 {0}(75,287)(25,287)(25,289)(17,289){1}
wire w17;    //: /sn:0 {0}(517,388)(479,388)(479,421)(249,421)(249,427){1}
//: {2}(247,429)(239,429){3}
//: {4}(249,431)(249,493)(62,493)(62,515)(77,515){5}
wire w12;    //: /sn:0 {0}(118,354)(142,354)(142,353)(194,353){1}
wire w11;    //: /sn:0 {0}(517,368)(469,368)(469,276)(246,276){1}
//: {2}(242,276)(234,276){3}
//: {4}(244,278)(244,332)(61,332)(61,345)(76,345){5}
wire w2;    //: /sn:0 {0}(517,338)(503,338)(503,41)(247,41){1}
//: {2}(243,41)(235,41){3}
//: {4}(245,43)(245,93)(65,93)(65,110)(80,110){5}
wire w5;    //: /sn:0 {0}(517,348)(492,348)(492,122)(247,122){1}
//: {2}(243,122)(235,122){3}
//: {4}(245,124)(245,174)(69,174)(69,193)(79,193){5}
wire w9;    //: /sn:0 {0}(117,277)(149,277)(149,276)(192,276){1}
wire w26;    //: /sn:0 {0}(80,129)(25,129)(25,126)(17,126){1}
//: enddecls

  MUX2 g8 (.in0(w25), .in1(w23), .c(ctrl), .out(w0));   //: @(81, 23) /sz:(40, 42) /sn:0 /p:[ Li0>1 Li1>0 Bi0>15 Ro0<0 ]
  FFD g4 (.D(w12), .Clk(clk), .Y(w14));   //: @(195, 334) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>23 Ro0<3 ]
  //: joint g51 (w17) @(249, 429) /w:[ -1 1 2 4 ]
  assign w36 = in[1]; //: TAP g37 @(11,533) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  assign w30 = in[4]; //: TAP g34 @(11,289) /sn:0 /R:2 /w:[ 1 9 10 ] /ss:1
  MUX2 g13 (.in0(w11), .in1(w32), .c(ctrl), .out(w12));   //: @(77, 336) /sz:(40, 42) /sn:0 /p:[ Li0>5 Li1>0 Bi0>23 Ro0<0 ]
  FFD g3 (.D(w9), .Clk(clk), .Y(w11));   //: @(193, 257) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>21 Ro0<3 ]
  FFD g2 (.D(w6), .Clk(clk), .Y(w8));   //: @(192, 184) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>19 Ro0<3 ]
  FFD g1 (.D(w7), .Clk(clk), .Y(w5));   //: @(194, 103) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>17 Ro0<3 ]
  //: OUT g16 (out) @(288,640) /sn:0 /w:[ 0 ]
  MUX2 g11 (.in0(w5), .in1(w28), .c(ctrl), .out(w6));   //: @(80, 184) /sz:(40, 42) /sn:0 /p:[ Li0>5 Li1>0 Bi0>19 Ro0<0 ]
  //: joint g50 (w1) @(242, 523) /w:[ -1 2 4 1 ]
  //: joint g28 (ctrl) @(375, 320) /w:[ -1 10 20 9 ]
  MUX2 g10 (.in0(w2), .in1(w26), .c(ctrl), .out(w7));   //: @(81, 101) /sz:(40, 42) /sn:0 /p:[ Li0>5 Li1>0 Bi0>17 Ro0<0 ]
  assign w26 = in[6]; //: TAP g32 @(11,126) /sn:0 /R:2 /w:[ 1 13 14 ] /ss:1
  //: joint g27 (ctrl) @(375, 389) /w:[ -1 8 22 7 ]
  //: joint g19 (clk) @(326, 395) /w:[ -1 8 22 7 ]
  FFD g38 (.D(w4), .Clk(clk), .Y(out));   //: @(194, 596) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>0 Ro0<5 ]
  FFD g6 (.D(w18), .Clk(clk), .Y(w1));   //: @(191, 504) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>27 Ro0<5 ]
  //: IN g7 (in) @(13,15) /sn:0 /R:3 /w:[ 17 ]
  //: GROUND g9 (w25) @(44,32) /sn:0 /R:3 /w:[ 0 ]
  assign w23 = in[7]; //: TAP g31 @(11,44) /sn:0 /R:2 /w:[ 1 15 16 ] /ss:1
  //: joint g20 (clk) @(326, 314) /w:[ -1 10 20 9 ]
  MUX2 g15 (.in0(w17), .in1(w36), .c(ctrl), .out(w18));   //: @(78, 506) /sz:(40, 42) /sn:0 /p:[ Li0>5 Li1>0 Bi0>27 Ro0<0 ]
  MUX2 g39 (.in0(w1), .in1(w16), .c(ctrl), .out(w4));   //: @(77, 594) /sz:(40, 42) /sn:0 /p:[ Li0>0 Li1>0 Bi0>0 Ro0<1 ]
  //: joint g48 (w14) @(246, 353) /w:[ 1 -1 2 4 ]
  assign putM = {w2, w5, w8, w11, w14, w17, w1, out}; //: CONCAT g43  @(522,373) /sn:0 /w:[ 1 0 0 0 0 0 0 3 3 ] /dr:0 /tp:0 /drp:1
  //: joint g29 (ctrl) @(375, 236) /w:[ -1 12 18 11 ]
  //: joint g25 (ctrl) @(375, 482) /w:[ -1 6 24 5 ]
  //: IN g17 (clk) @(326,689) /sn:0 /R:1 /w:[ 29 ]
  //: OUT g52 (putM) @(599,380) /sn:0 /w:[ 0 ]
  assign w16 = in[0]; //: TAP g42 @(11,622) /sn:0 /R:2 /anc:1 /w:[ 1 1 2 ] /ss:1
  MUX2 g14 (.in0(w14), .in1(w34), .c(ctrl), .out(w15));   //: @(76, 410) /sz:(40, 42) /sn:0 /p:[ Li0>5 Li1>0 Bi0>25 Ro0<0 ]
  FFD g5 (.D(w15), .Clk(clk), .Y(w17));   //: @(198, 410) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>25 Ro0<3 ]
  //: joint g47 (w11) @(244, 276) /w:[ 1 -1 2 4 ]
  //: joint g44 (w2) @(245, 41) /w:[ 1 -1 2 4 ]
  assign w34 = in[2]; //: TAP g36 @(11,437) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  //: joint g24 (clk) @(326, 560) /w:[ -1 4 26 3 ]
  //: joint g21 (clk) @(326, 242) /w:[ -1 12 18 11 ]
  //: joint g41 (ctrl) @(375, 656) /w:[ -1 2 1 28 ]
  //: IN g23 (ctrl) @(375,685) /sn:0 /R:1 /w:[ 29 ]
  //: joint g40 (clk) @(326, 667) /w:[ -1 2 1 28 ]
  //: joint g46 (w8) @(243, 203) /w:[ 1 -1 2 4 ]
  //: joint g45 (w5) @(245, 122) /w:[ 1 -1 2 4 ]
  assign w32 = in[3]; //: TAP g35 @(11,362) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  //: joint g26 (ctrl) @(375, 549) /w:[ -1 4 26 3 ]
  //: joint g22 (clk) @(326, 161) /w:[ -1 14 16 13 ]
  FFD g0 (.D(w0), .Clk(clk), .Y(w2));   //: @(194, 22) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>15 Ro0<3 ]
  //: joint g18 (clk) @(326, 469) /w:[ -1 6 24 5 ]
  MUX2 g12 (.in0(w8), .in1(w30), .c(ctrl), .out(w9));   //: @(76, 259) /sz:(40, 42) /sn:0 /p:[ Li0>5 Li1>0 Bi0>21 Ro0<0 ]
  assign w28 = in[5]; //: TAP g33 @(11,211) /sn:0 /R:2 /w:[ 1 11 12 ] /ss:1
  //: joint g30 (ctrl) @(375, 151) /w:[ -1 14 16 13 ]
  //: joint g49 (out) @(250, 618) /w:[ 2 4 -1 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFD
module FFD(Clk, Y, D);
//: interface  /sz:(40, 40) /bd:[ Li0>D(19/40) Bi0>Clk(18/40) Ro0<Y(19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Clk;    //: /sn:0 {0}(375,157)(404,157)(404,154)(414,154){1}
//: {2}(416,152)(416,137)(418,137)(418,124){3}
//: {4}(416,156)(416,189){5}
input D;    //: /sn:0 {0}(238,101)(278,101){1}
output Y;    //: /sn:0 {0}(441,102)(470,102)(470,101)(485,101){1}
wire w1;    //: /sn:0 {0}(333,158)(297,158)(297,123){1}
wire w2;    //: /sn:0 {0}(320,101)(384,101)(384,102)(399,102){1}
//: enddecls

  //: joint g4 (Clk) @(416, 154) /w:[ -1 2 1 4 ]
  INV1 g3 (.in(Clk), .out(w1));   //: @(334, 138) /sz:(40, 40) /R:2 /sn:0 /p:[ Ri0>0 Lo0<0 ]
  //: IN g2 (Clk) @(416,191) /sn:0 /R:1 /w:[ 5 ]
  FFDLS g1 (.D(w2), .Clk(Clk), .Y(Y));   //: @(400, 83) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>3 Ro0<0 ]
  //: OUT g6 (Y) @(482,101) /sn:0 /w:[ 1 ]
  //: IN g5 (D) @(236,101) /sn:0 /w:[ 0 ]
  FFDLS g0 (.D(D), .Clk(w1), .Y(w2));   //: @(279, 82) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin BySaddsub2
module BySaddsub2(S, load, B2, clk, B, A, A2, mode);
//: interface  /sz:(73, 80) /bd:[ Ti0>B[7:0](54/73) Ti1>A[7:0](12/73) Li0>clk(63/80) Li1>load(21/80) Ri0>mode(22/80) Bo0<S[8:0](37/73) Ro0<A2[7:0](50/80) Ro1<B2[7:0](74/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:565,126)(472,126)(472,157)(457,157){1}
input [7:0] A;    //: /sn:0 {0}(#:39,140)(106,140)(106,141)(#:121,141){1}
output [7:0] A2;    //: /sn:0 {0}(244,101)(187,101)(#:187,140)(172,140){1}
input mode;    //: /sn:0 {0}(678,272)(678,209)(678,209)(678,199){1}
//: {2}(680,197)(697,197){3}
//: {4}(676,197)(448,197){5}
//: {6}(444,197)(391,197)(391,413)(169,413)(169,336)(180,336){7}
//: {8}(446,199)(446,219)(417,219)(417,190){9}
output [7:0] B2;    //: /sn:0 {0}(#:478,236)(359,236)(359,190){1}
input load;    //: /sn:0 {0}(635,105)(635,76)(636,76)(636,67){1}
//: {2}(638,65)(688,65){3}
//: {4}(634,65)(448,65){5}
//: {6}(444,65)(87,65)(87,246){7}
//: {8}(89,248)(131,248)(131,175){9}
//: {10}(87,250)(87,375)(198,375)(198,351){11}
//: {12}(446,67)(446,109)(417,109)(417,132){13}
input clk;    //: /sn:0 {0}(478,432)(457,432)(457,386){1}
//: {2}(457,382)(457,296)(521,296)(521,40){3}
//: {4}(523,38)(687,38){5}
//: {6}(519,38)(409,38){7}
//: {8}(405,38)(146,38)(146,91){9}
//: {10}(407,40)(407,80)(378,80)(378,132){11}
//: {12}(455,384)(342,384)(342,362){13}
output [8:0] S;    //: /sn:0 {0}(#:598,433)(564,433)(564,378)(#:539,378){1}
wire w14;    //: /sn:0 {0}(524,361)(524,329)(679,329)(679,314){1}
wire w3;    //: /sn:0 {0}(163,175)(163,198)(278,198)(278,213){1}
wire w0;    //: /sn:0 {0}(613,291)(613,310)(490,310)(490,361){1}
wire w1;    //: /sn:0 {0}(641,147)(641,234)(622,234)(622,249){1}
wire w8;    //: /sn:0 {0}(338,157)(305,157)(305,213){1}
wire w2;    //: /sn:0 {0}(602,249)(602,239)(534,239)(534,286)(297,286)(297,271){1}
wire w12;    //: /sn:0 {0}(271,243)(165,243)(165,317)(180,317){1}
wire w11;    //: /sn:0 {0}(318,247)(372,247)(372,340)(365,340){1}
wire w9;    //: /sn:0 {0}(222,326)(258,326)(258,340)(323,340){1}
//: enddecls

  //: joint g8 (clk) @(521, 38) /w:[ 4 -1 6 3 ]
  MUX2 g4 (.in0(w12), .in1(mode), .c(load), .out(w9));   //: @(181, 308) /sz:(40, 42) /sn:0 /p:[ Li0>1 Li1>7 Bi0>11 Ro0<0 ]
  //: joint g13 (mode) @(446, 197) /w:[ 5 -1 6 8 ]
  FFD g3 (.D(w9), .Clk(clk), .Y(w11));   //: @(324, 321) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>13 Ro0<1 ]
  FA g2 (.A(w3), .B(w8), .Cin(w11), .Cout(w12), .S(w2));   //: @(272, 214) /sz:(45, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<1 ]
  REG8sINaddsub g1 (.clk(clk), .ctrl(load), .mode(mode), .in(B), .out(w8), .Out2(B2));   //: @(340, 133) /sz:(117, 56) /R:3 /sn:0 /p:[ Ti0>11 Ti1>13 Bi0>9 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g11 (load) @(87, 248) /w:[ 8 7 -1 10 ]
  //: OUT g16 (S) @(595,433) /sn:0 /w:[ 0 ]
  //: IN g10 (load) @(690,65) /sn:0 /R:2 /w:[ 3 ]
  //: OUT g19 (B2) @(475,236) /sn:0 /w:[ 0 ]
  //: IN g6 (clk) @(689,38) /sn:0 /R:2 /w:[ 5 ]
  //: joint g7 (clk) @(407, 38) /w:[ 7 -1 8 10 ]
  //: joint g9 (clk) @(457, 384) /w:[ -1 2 12 1 ]
  //: joint g20 (load) @(636, 65) /w:[ 2 -1 4 1 ]
  //: IN g15 (B) @(567,126) /sn:0 /R:2 /w:[ 0 ]
  //: joint g17 (load) @(446, 65) /w:[ 5 -1 6 12 ]
  //: IN g14 (A) @(37,140) /sn:0 /w:[ 0 ]
  REG9sOUT g5 (.ctrlNeg(w14), .in(w0), .clk(clk), .out(S));   //: @(479, 362) /sz:(59, 90) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>0 Ro0<1 ]
  INV1 g21 (.in(load), .out(w1));   //: @(616, 106) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  INV1 g24 (.in(mode), .out(w14));   //: @(659, 273) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  //: joint g23 (mode) @(678, 197) /w:[ 2 -1 4 1 ]
  AND2 g22 (.in1(w1), .in2(w2), .out(w0));   //: @(592, 250) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<0 ]
  REG8sIN g0 (.clk(clk), .in(A), .ctrl(load), .out(w3), .putM(A2));   //: @(122, 92) /sz:(49, 82) /sn:0 /p:[ Ti0>9 Li0>1 Bi0>9 Bo0<0 Ro0<1 ]
  //: OUT g18 (A2) @(241,101) /sn:0 /w:[ 0 ]
  //: IN g12 (mode) @(699,197) /sn:0 /R:2 /w:[ 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux8
module Mux8(A1, B, B2, A, ctrl);
//: interface  /sz:(63, 80) /bd:[ Ti0>ctrl(32/63) Li0>A[7:0](16/80) Li1>B[7:0](64/80) Ro0<A1[7:0](16/80) Ro1<B2[7:0](64/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:1047,108)(1030,108){1}
//: {2}(1029,108)(967,108){3}
//: {4}(966,108)(911,108){5}
//: {6}(910,108)(860,108){7}
//: {8}(859,108)(803,108){9}
//: {10}(802,108)(754,108){11}
//: {12}(753,108)(698,108){13}
//: {14}(697,108)(639,108){15}
//: {16}(638,108)(#:583,108){17}
supply0 w56;    //: /sn:0 {0}(949,354)(949,237)(940,237)(940,140){1}
//: {2}(942,138)(997,138){3}
//: {4}(1001,138)(1034,138){5}
//: {6}(999,140)(999,150)(1012,150)(1012,382){7}
//: {8}(938,138)(884,138){9}
//: {10}(880,138)(827,138){11}
//: {12}(823,138)(778,138){13}
//: {14}(774,138)(724,138){15}
//: {16}(720,138)(678,138){17}
//: {18}(674,138)(614,138){19}
//: {20}(610,138)(533,138){21}
//: {22}(529,138)(478,138){23}
//: {24}(474,138)(422,138){25}
//: {26}(418,138)(368,138){27}
//: {28}(364,138)(318,138){29}
//: {30}(314,138)(264,138){31}
//: {32}(260,138)(209,138){33}
//: {34}(205,138)(150,138){35}
//: {36}(146,138)(56,138){37}
//: {38}(148,140)(148,150)(156,150)(156,165){39}
//: {40}(207,140)(207,150)(218,150)(218,199){41}
//: {42}(262,140)(262,150)(278,150)(278,232){43}
//: {44}(316,140)(316,150)(332,150)(332,260){45}
//: {46}(366,140)(366,150)(382,150)(382,296){47}
//: {48}(420,140)(420,150)(444,150)(444,327){49}
//: {50}(476,140)(476,150)(497,150)(497,356){51}
//: {52}(531,140)(531,150)(550,150)(550,379){53}
//: {54}(612,140)(612,150)(621,150)(621,160){55}
//: {56}(676,140)(676,150)(680,150)(680,183){57}
//: {58}(722,140)(722,150)(734,150)(734,219){59}
//: {60}(776,140)(776,150)(786,150)(786,250){61}
//: {62}(825,140)(825,150)(841,150)(841,285){63}
//: {64}(882,140)(882,150)(891,150)(891,323){65}
input [7:0] A;    //: /sn:0 {0}(#:103,125)(173,125){1}
//: {2}(174,125)(236,125){3}
//: {4}(237,125)(295,125){5}
//: {6}(296,125)(349,125){7}
//: {8}(350,125)(399,125){9}
//: {10}(400,125)(461,125){11}
//: {12}(462,125)(514,125){13}
//: {14}(515,125)(567,125){15}
//: {16}(568,125)(601,125){17}
output [7:0] B2;    //: /sn:0 {0}(734,581)(842,581)(#:842,573){1}
input ctrl;    //: /sn:0 {0}(27,47)(65,47)(65,63){1}
output [7:0] A1;    //: /sn:0 {0}(266,539)(349,539)(#:349,522){1}
wire w6;    //: /sn:0 {0}(640,160)(640,120)(639,120)(639,112){1}
wire w7;    //: /sn:0 {0}(228,241)(228,490)(324,490)(324,516){1}
wire w45;    //: /sn:0 {0}(910,323)(910,120)(911,120)(911,112){1}
wire w14;    //: /sn:0 {0}(631,202)(631,552)(807,552)(807,567){1}
wire w15;    //: /sn:0 {0}(344,516)(344,432)(342,432)(342,302){1}
wire w19;    //: /sn:0 {0}(354,516)(354,434)(392,434)(392,338){1}
wire w51;    //: /sn:0 {0}(867,567)(867,505)(959,505)(959,396){1}
wire w0;    //: /sn:0 {0}(66,105)(66,182){1}
//: {2}(68,184)(606,184){3}
//: {4}(64,184)(42,184)(42,222)(93,222){5}
//: {6}(97,222)(107,222)(107,223)(203,223){7}
//: {8}(95,220)(95,188)(107,188)(107,189)(141,189){9}
//: {10}(95,224)(95,255){11}
//: {12}(97,257)(107,257)(107,256)(263,256){13}
//: {14}(97,257)(87,257)(87,207)(665,207){15}
//: {16}(95,259)(95,281){17}
//: {18}(97,283)(107,283)(107,284)(317,284){19}
//: {20}(97,283)(87,283)(87,243)(719,243){21}
//: {22}(95,285)(95,318){23}
//: {24}(97,320)(367,320){25}
//: {26}(97,320)(87,320)(87,274)(771,274){27}
//: {28}(95,322)(95,349){29}
//: {30}(97,351)(429,351){31}
//: {32}(97,351)(87,351)(87,309)(826,309){33}
//: {34}(95,353)(95,377){35}
//: {36}(97,379)(107,379)(107,380)(482,380){37}
//: {38}(97,379)(87,379)(87,347)(876,347){39}
//: {40}(95,381)(95,399){41}
//: {42}(97,401)(107,401)(107,403)(535,403){43}
//: {44}(97,401)(87,401)(87,378)(934,378){45}
//: {46}(95,403)(95,434)(107,434)(107,406)(997,406){47}
wire w3;    //: /sn:0 {0}(166,207)(166,501)(314,501)(314,516){1}
wire w37;    //: /sn:0 {0}(805,250)(805,120)(803,120)(803,112){1}
wire w21;    //: /sn:0 {0}(463,327)(463,137)(462,137)(462,129){1}
wire w43;    //: /sn:0 {0}(847,567)(847,491)(851,491)(851,327){1}
wire w31;    //: /sn:0 {0}(384,516)(384,491)(560,491)(560,421){1}
wire w23;    //: /sn:0 {0}(364,516)(364,450)(454,450)(454,369){1}
wire w41;    //: /sn:0 {0}(860,285)(860,112){1}
wire w1;    //: /sn:0 {0}(175,165)(175,137)(174,137)(174,129){1}
wire w25;    //: /sn:0 {0}(516,356)(516,137)(515,137)(515,129){1}
wire w35;    //: /sn:0 {0}(744,261)(744,535)(827,535)(827,567){1}
wire w30;    //: /sn:0 {0}(690,225)(690,546)(817,546)(817,567){1}
wire w17;    //: /sn:0 {0}(401,296)(401,137)(400,137)(400,129){1}
wire w22;    //: /sn:0 {0}(699,183)(699,120)(698,120)(698,112){1}
wire w53;    //: /sn:0 {0}(1031,382)(1031,120)(1030,120)(1030,112){1}
wire w11;    //: /sn:0 {0}(288,274)(288,481)(334,481)(334,516){1}
wire w49;    //: /sn:0 {0}(968,354)(968,120)(967,120)(967,112){1}
wire w13;    //: /sn:0 {0}(351,260)(351,137)(350,137)(350,129){1}
wire w27;    //: /sn:0 {0}(374,516)(374,465)(507,465)(507,398){1}
wire w5;    //: /sn:0 {0}(237,199)(237,129){1}
wire w33;    //: /sn:0 {0}(753,219)(753,120)(754,120)(754,112){1}
wire w29;    //: /sn:0 {0}(569,379)(569,137)(568,137)(568,129){1}
wire w47;    //: /sn:0 {0}(857,567)(857,491)(901,491)(901,365){1}
wire w9;    //: /sn:0 {0}(297,232)(297,137)(296,137)(296,129){1}
wire w39;    //: /sn:0 {0}(837,567)(837,482)(796,482)(796,292){1}
wire w55;    //: /sn:0 {0}(877,567)(877,528)(1022,528)(1022,424){1}
//: enddecls

  MUX2 g4 (.in0(w9), .in1(w56), .c(w0), .out(w11));   //: @(264, 233) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>43 Li0>13 Bo0<0 ]
  MUX2 g8 (.in0(w25), .in1(w56), .c(w0), .out(w27));   //: @(483, 357) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>51 Li0>37 Bo0<1 ]
  //: OUT g61 (A1) @(269,539) /sn:0 /R:2 /w:[ 0 ]
  MUX2 g3 (.in0(w5), .in1(w56), .c(w0), .out(w7));   //: @(204, 200) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>41 Li0>7 Bo0<0 ]
  assign w13 = A[3]; //: TAP g13 @(350,123) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  MUX2 g34 (.in0(w53), .in1(w56), .c(w0), .out(w55));   //: @(998, 383) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>7 Li0>47 Bo0<1 ]
  assign w33 = B[2]; //: TAP g37 @(754,106) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  //: joint g51 (w56) @(612, 138) /w:[ 19 -1 20 54 ]
  //: joint g55 (w56) @(776, 138) /w:[ 13 -1 14 60 ]
  //: joint g58 (w56) @(940, 138) /w:[ 2 -1 8 1 ]
  MUX2 g2 (.in0(w1), .in1(w56), .c(w0), .out(w3));   //: @(142, 166) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>39 Li0>9 Bo0<0 ]
  //: joint g59 (w56) @(999, 138) /w:[ 4 -1 3 6 ]
  //: IN g1 (B) @(581,108) /sn:0 /w:[ 17 ]
  //: joint g64 (w0) @(66, 184) /w:[ 2 1 4 -1 ]
  assign w5 = A[1]; //: TAP g11 @(237,123) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w25 = A[6]; //: TAP g16 @(515,123) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  assign w1 = A[0]; //: TAP g10 @(174,123) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  MUX2 g28 (.in0(w22), .in1(w56), .c(w0), .out(w30));   //: @(666, 184) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>57 Li0>15 Bo0<0 ]
  //: joint g50 (w56) @(476, 138) /w:[ 23 -1 24 50 ]
  //: joint g19 (w0) @(95, 401) /w:[ 42 41 44 46 ]
  MUX2 g27 (.in0(w6), .in1(w56), .c(w0), .out(w14));   //: @(607, 161) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>55 Li0>3 Bo0<0 ]
  MUX2 g32 (.in0(w45), .in1(w56), .c(w0), .out(w47));   //: @(877, 324) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>65 Li0>39 Bo0<1 ]
  MUX2 g6 (.in0(w17), .in1(w56), .c(w0), .out(w19));   //: @(368, 297) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>47 Li0>25 Bo0<1 ]
  assign w37 = B[3]; //: TAP g38 @(803,106) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  MUX2 g7 (.in0(w21), .in1(w56), .c(w0), .out(w23));   //: @(430, 328) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>49 Li0>31 Bo0<1 ]
  MUX2 g9 (.in0(w29), .in1(w56), .c(w0), .out(w31));   //: @(536, 380) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>53 Li0>43 Bo0<1 ]
  //: joint g53 (w56) @(531, 138) /w:[ 21 -1 22 52 ]
  //: joint g57 (w56) @(882, 138) /w:[ 9 -1 10 64 ]
  assign w21 = A[5]; //: TAP g15 @(462,123) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  //: joint g20 (w0) @(95, 379) /w:[ 36 35 38 40 ]
  MUX2 g31 (.in0(w41), .in1(w56), .c(w0), .out(w43));   //: @(827, 286) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>63 Li0>33 Bo0<1 ]
  assign w41 = B[4]; //: TAP g39 @(860,106) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: GROUND g43 (w56) @(50,138) /sn:0 /R:3 /w:[ 37 ]
  //: joint g48 (w56) @(366, 138) /w:[ 27 -1 28 46 ]
  assign w29 = A[7]; //: TAP g17 @(568,123) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  //: joint g25 (w0) @(95, 222) /w:[ 6 8 5 10 ]
  MUX2 g29 (.in0(w33), .in1(w56), .c(w0), .out(w35));   //: @(720, 220) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>59 Li0>21 Bo0<0 ]
  assign B2 = {w55, w51, w47, w43, w39, w35, w30, w14}; //: CONCAT g62  @(842,572) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 1 1 1 ] /dr:0 /tp:0 /drp:1
  assign w53 = B[7]; //: TAP g42 @(1030,106) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: joint g52 (w56) @(676, 138) /w:[ 17 -1 18 56 ]
  //: OUT g63 (B2) @(737,581) /sn:0 /R:2 /w:[ 0 ]
  MUX2 g5 (.in0(w13), .in1(w56), .c(w0), .out(w15));   //: @(318, 261) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>45 Li0>19 Bo0<1 ]
  assign w17 = A[4]; //: TAP g14 @(400,123) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  //: joint g56 (w56) @(825, 138) /w:[ 11 -1 12 62 ]
  //: joint g44 (w56) @(148, 138) /w:[ 35 -1 36 38 ]
  //: joint g47 (w56) @(316, 138) /w:[ 29 -1 30 44 ]
  //: joint g21 (w0) @(95, 351) /w:[ 30 29 32 34 ]
  //: joint g24 (w0) @(95, 257) /w:[ 12 11 14 16 ]
  assign w22 = B[1]; //: TAP g36 @(698,106) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  //: joint g23 (w0) @(95, 283) /w:[ 18 17 20 22 ]
  assign w49 = B[6]; //: TAP g41 @(967,106) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  assign w45 = B[5]; //: TAP g40 @(911,106) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: joint g54 (w56) @(722, 138) /w:[ 15 -1 16 58 ]
  assign A1 = {w31, w27, w23, w19, w15, w11, w7, w3}; //: CONCAT g60  @(349,521) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 1 1 1 ] /dr:0 /tp:0 /drp:1
  INV1 g26 (.in(ctrl), .out(w0));   //: @(46, 64) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>1 Bo0<0 ]
  //: IN g0 (A) @(101,125) /sn:0 /w:[ 0 ]
  //: joint g22 (w0) @(95, 320) /w:[ 24 23 26 28 ]
  assign w6 = B[0]; //: TAP g35 @(639,106) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  //: joint g45 (w56) @(207, 138) /w:[ 33 -1 34 40 ]
  //: joint g46 (w56) @(262, 138) /w:[ 31 -1 32 42 ]
  assign w9 = A[2]; //: TAP g12 @(296,123) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: IN g18 (ctrl) @(25,47) /sn:0 /w:[ 0 ]
  MUX2 g30 (.in0(w37), .in1(w56), .c(w0), .out(w39));   //: @(772, 251) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>61 Li0>27 Bo0<1 ]
  MUX2 g33 (.in0(w49), .in1(w56), .c(w0), .out(w51));   //: @(935, 355) /sz:(42, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>45 Bo0<1 ]
  //: joint g49 (w56) @(420, 138) /w:[ 25 -1 26 48 ]

endmodule
//: /netlistEnd

//: /netlistBegin LATCHSR
module LATCHSR(Y1, r, s, Y);
//: interface  /sz:(81, 47) /bd:[ Li0>s(7/47) Li1>r(31/47) Ro0<Y1(10/47) Ro1<Y(31/47) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input r;    //: /sn:0 {0}(253,213)(211,213)(211,215)(196,215){1}
input s;    //: /sn:0 {0}(255,113)(214,113)(214,111)(199,111){1}
output Y1;    //: /sn:0 {0}(297,123)(305,123){1}
//: {2}(309,123)(350,123)(350,121)(389,121){3}
//: {4}(307,125)(307,167)(238,167)(238,191)(253,191){5}
output Y;    //: /sn:0 {0}(255,135)(245,135)(245,148)(318,148)(318,199){1}
//: {2}(320,201)(330,201)(330,193)(380,193){3}
//: {4}(316,201)(295,201){5}
//: enddecls

  //: OUT g4 (Y1) @(386,121) /sn:0 /w:[ 3 ]
  //: IN g3 (r) @(194,215) /sn:0 /w:[ 1 ]
  //: IN g2 (s) @(197,111) /sn:0 /w:[ 1 ]
  NOR2 g1 (.in2(r), .in1(Y1), .out(Y));   //: @(254, 183) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>5 Ro0<5 ]
  //: joint g6 (Y) @(318, 201) /w:[ 2 1 4 -1 ]
  //: joint g7 (Y1) @(307, 123) /w:[ 2 -1 1 4 ]
  //: OUT g5 (Y) @(377,193) /sn:0 /w:[ 3 ]
  NOR2 g0 (.in2(Y), .in1(s), .out(Y1));   //: @(256, 105) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin NOR2
module NOR2(in1, out, in2);
//: interface  /sz:(40, 40) /bd:[ Li0>in2(30/40) Li1>in1(8/40) Ro0<out(18/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output out;    //: /sn:0 {0}(269,219)(269,227)(269,227)(269,235){1}
//: {2}(267,237)(187,237)(187,237)(343,237){3}
//: {4}(269,239)(269,261)(269,261)(269,269){5}
//: {6}(271,271)(332,271)(332,286){7}
//: {8}(267,271)(235,271)(235,302){9}
supply1 w0;    //: /sn:0 {0}(269,97)(269,122)(269,122)(269,137){1}
supply0 w1;    //: /sn:0 {0}(270,365)(270,343)(270,343)(270,333){1}
//: {2}(272,331)(332,331)(332,303){3}
//: {4}(268,331)(235,331)(235,319){5}
input in1;    //: /sn:0 {0}(144,145)(176,145)(176,145)(189,145){1}
//: {2}(193,145)(242,145)(242,145)(255,145){3}
//: {4}(191,147)(191,294)(318,294){5}
input in2;    //: /sn:0 {0}(142,210)(162,210)(162,210)(157,210){1}
//: {2}(161,210)(207,210)(207,210)(255,210){3}
//: {4}(159,212)(159,310)(221,310){5}
wire w2;    //: /sn:0 {0}(269,154)(269,187)(269,187)(269,202){1}
//: enddecls

  _GGNMOS #(2, 1) g4 (.Z(out), .S(w1), .G(in2));   //: @(229,310) /sn:0 /w:[ 9 5 5 ]
  //: IN g8 (in1) @(142,145) /sn:0 /w:[ 0 ]
  _GGPMOS #(2, 1) g3 (.Z(out), .S(w2), .G(in2));   //: @(263,210) /sn:0 /w:[ 0 1 3 ]
  //: joint g13 (in2) @(159, 210) /w:[ 2 -1 1 4 ]
  _GGPMOS #(2, 1) g2 (.Z(w2), .S(w0), .G(in1));   //: @(263,145) /sn:0 /w:[ 0 1 3 ]
  //: GROUND g1 (w1) @(270,371) /sn:0 /w:[ 0 ]
  //: joint g11 (out) @(269, 237) /w:[ -1 1 2 4 ]
  //: OUT g10 (out) @(340,237) /sn:0 /w:[ 3 ]
  //: joint g6 (w1) @(270, 331) /w:[ 2 -1 4 1 ]
  //: joint g7 (out) @(269, 271) /w:[ 6 5 8 -1 ]
  //: IN g9 (in2) @(140,210) /sn:0 /w:[ 0 ]
  _GGNMOS #(2, 1) g5 (.Z(out), .S(w1), .G(in1));   //: @(326,294) /sn:0 /w:[ 7 3 5 ]
  //: VDD g0 (w0) @(280,97) /sn:0 /w:[ 0 ]
  //: joint g12 (in1) @(191, 145) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFDLS
module FFDLS(Clk, D, Y);
//: interface  /sz:(40, 40) /bd:[ Li0>D(19/40) Bi0>Clk(18/40) Ro0<Y(19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Clk;    //: /sn:0 {0}(380,218)(405,218)(405,158){1}
input D;    //: /sn:0 {0}(268,145)(215,145)(215,116){1}
//: {2}(217,114)(374,114)(374,124)(387,124){3}
//: {4}(213,114)(172,114){5}
output Y;    //: /sn:0 {0}(523,139)(444,139)(444,135)(429,135){1}
wire w0;    //: /sn:0 {0}(387,145)(325,145)(325,144)(310,144){1}
//: enddecls

  //: IN g4 (Clk) @(378,218) /sn:0 /w:[ 0 ]
  //: joint g3 (D) @(215, 114) /w:[ 2 -1 4 1 ]
  //: IN g2 (D) @(170,114) /sn:0 /w:[ 5 ]
  INV1 g1 (.in(D), .out(w0));   //: @(269, 124) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  //: OUT g5 (Y) @(520,139) /sn:0 /w:[ 0 ]
  FFSR g0 (.S(D), .R(w0), .clk(Clk), .Y(Y));   //: @(388, 117) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>0 Bi0>1 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA
module FA(Cin, S, Cout, B, A);
//: interface  /sz:(45, 56) /bd:[ Ti0>B(33/45) Ti1>A(6/45) Ri0>Cin(33/56) Lo0<Cout(29/56) Bo0<S(25/45) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(168,243)(120,243)(120,154){1}
//: {2}(122,152)(171,152)(171,138)(184,138){3}
//: {4}(118,152)(92,152){5}
input A;    //: /sn:0 {0}(95,110)(150,110){1}
//: {2}(154,110)(173,110)(173,120)(184,120){3}
//: {4}(152,112)(152,223)(168,223){5}
output Cout;    //: /sn:0 {0}(442,254)(381,254){1}
input Cin;    //: /sn:0 {0}(280,324)(263,324)(263,192){1}
//: {2}(265,190)(308,190)(308,152)(321,152){3}
//: {4}(261,190)(92,190){5}
output S;    //: /sn:0 {0}(448,152)(413,152)(413,151)(378,151){1}
wire w6;    //: /sn:0 {0}(322,332)(329,332)(329,266)(339,266){1}
wire w3;    //: /sn:0 {0}(210,231)(324,231)(324,246)(339,246){1}
wire w2;    //: /sn:0 {0}(280,344)(271,344)(271,139){1}
//: {2}(273,137)(308,137)(308,134)(321,134){3}
//: {4}(269,137)(241,137){5}
//: enddecls

  NAND2 g8 (.in2(w2), .in1(Cin), .out(w6));   //: @(281, 314) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  //: IN g4 (Cin) @(90,190) /sn:0 /w:[ 5 ]
  //: OUT g3 (S) @(445,152) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(120, 152) /w:[ 2 -1 4 1 ]
  //: OUT g2 (Cout) @(439,254) /sn:0 /w:[ 0 ]
  //: IN g1 (B) @(90,152) /sn:0 /w:[ 5 ]
  //: joint g11 (w2) @(271, 137) /w:[ 2 -1 4 1 ]
  //: joint g10 (Cin) @(263, 190) /w:[ 2 -1 4 1 ]
  EXOR2 g6 (.a(w2), .b(Cin), .out(S));   //: @(322, 124) /sz:(55, 42) /sn:0 /p:[ Li0>3 Li1>3 Ro0<1 ]
  NAND2 g9 (.in2(w6), .in1(w3), .out(Cout));   //: @(340, 236) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 ]
  NAND2 g7 (.in2(B), .in1(A), .out(w3));   //: @(169, 213) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>5 Ro0<0 ]
  EXOR2 g5 (.a(A), .b(B), .out(w2));   //: @(185, 110) /sz:(55, 42) /sn:0 /p:[ Li0>3 Li1>3 Ro0<5 ]
  //: IN g0 (A) @(93,110) /sn:0 /w:[ 0 ]
  //: joint g12 (A) @(152, 110) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin REG9sOUT
module REG9sOUT(in, clk, out, ctrlNeg);
//: interface  /sz:(59, 90) /bd:[ Ti0>ctrlNeg(45/59) Ti1>in(11/59) Li0>clk(70/90) Ro0<out[8:0](16/90) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input in;    //: /sn:0 {0}(78,67)(157,67)(157,69)(172,69){1}
output [8:0] out;    //: /sn:0 {0}(#:432,385)(475,385)(475,335)(485,335){1}
input clk;    //: /sn:0 {0}(189,749)(189,759)(39,759)(39,675){1}
//: {2}(41,673)(188,673)(188,658){3}
//: {4}(39,671)(39,595){5}
//: {6}(41,593)(189,593)(189,584){7}
//: {8}(39,591)(39,526){9}
//: {10}(41,524)(188,524)(188,509){11}
//: {12}(39,522)(39,450){13}
//: {14}(41,448)(188,448)(188,431){15}
//: {16}(39,446)(39,368){17}
//: {18}(41,366)(190,366)(190,351){19}
//: {20}(39,364)(39,277){21}
//: {22}(41,275)(189,275)(189,262){23}
//: {24}(39,273)(39,190){25}
//: {26}(41,188)(190,188)(190,175){27}
//: {28}(39,186)(39,111){29}
//: {30}(41,109)(191,109)(191,91){31}
//: {32}(39,107)(39,80){33}
input ctrlNeg;    //: /sn:0 {0}(588,69)(425,69)(425,107){1}
wire w6;    //: /sn:0 {0}(169,487)(160,487)(160,459)(258,459)(258,411){1}
//: {2}(260,409)(274,409)(274,385)(426,385){3}
//: {4}(256,409)(211,409){5}
wire w7;    //: /sn:0 {0}(170,240)(163,240)(163,203)(264,203)(264,155){1}
//: {2}(266,153)(407,153)(407,355)(426,355){3}
//: {4}(262,153)(213,153){5}
wire w4;    //: /sn:0 {0}(170,562)(163,562)(163,535)(265,535)(265,489){1}
//: {2}(267,487)(315,487)(315,395)(426,395){3}
//: {4}(263,487)(211,487){5}
wire w0;    //: /sn:0 {0}(212,727)(417,727)(417,425)(426,425){1}
wire w3;    //: /sn:0 {0}(169,636)(159,636)(159,604)(258,604)(258,564){1}
//: {2}(260,562)(349,562)(349,405)(426,405){3}
//: {4}(256,562)(212,562){5}
wire w1;    //: /sn:0 {0}(170,727)(160,727)(160,695)(258,695)(258,638){1}
//: {2}(260,636)(408,636)(408,415)(426,415){3}
//: {4}(256,636)(211,636){5}
wire w8;    //: /sn:0 {0}(416,149)(416,345)(426,345){1}
wire w2;    //: /sn:0 {0}(405,107)(405,69)(264,69){1}
//: {2}(260,69)(214,69){3}
//: {4}(262,71)(262,122)(162,122)(162,153)(171,153){5}
wire w10;    //: /sn:0 {0}(169,409)(163,409)(163,379)(259,379)(259,331){1}
//: {2}(261,329)(387,329)(387,375)(426,375){3}
//: {4}(257,329)(213,329){5}
wire w9;    //: /sn:0 {0}(171,329)(162,329)(162,289)(256,289)(256,242){1}
//: {2}(258,240)(397,240)(397,365)(426,365){3}
//: {4}(254,240)(212,240){5}
//: enddecls

  //: IN g8 (in) @(76,67) /sn:0 /w:[ 0 ]
  FFD g4 (.D(w10), .Clk(clk), .Y(w6));   //: @(170, 390) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>15 Ro0<5 ]
  //: joint g13 (w10) @(259, 329) /w:[ 2 -1 4 1 ]
  FFD g3 (.D(w9), .Clk(clk), .Y(w10));   //: @(172, 310) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>19 Ro0<5 ]
  FFD g2 (.D(w7), .Clk(clk), .Y(w9));   //: @(171, 221) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>23 Ro0<5 ]
  FFD g1 (.D(w2), .Clk(clk), .Y(w7));   //: @(172, 134) /sz:(40, 40) /sn:0 /p:[ Li0>5 Bi0>27 Ro0<5 ]
  //: joint g16 (w3) @(258, 562) /w:[ 2 -1 4 1 ]
  //: joint g11 (w7) @(264, 153) /w:[ 2 -1 4 1 ]
  //: joint g28 (clk) @(39, 275) /w:[ 22 24 -1 21 ]
  AND2 g10 (.in2(w2), .in1(ctrlNeg), .out(w8));   //: @(395, 108) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<0 ]
  //: joint g19 (clk) @(39, 673) /w:[ 2 4 -1 1 ]
  //: joint g32 (clk) @(39, 593) /w:[ 6 8 -1 5 ]
  //: joint g27 (clk) @(39, 188) /w:[ 26 28 -1 25 ]
  FFD g6 (.D(w4), .Clk(clk), .Y(w3));   //: @(171, 543) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>7 Ro0<5 ]
  FFD g7 (.D(w3), .Clk(clk), .Y(w1));   //: @(170, 617) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>3 Ro0<5 ]
  assign out = {w8, w7, w9, w10, w6, w4, w3, w1, w0}; //: CONCAT g9  @(431,385) /sn:0 /w:[ 0 1 3 3 3 3 3 3 3 1 ] /dr:0 /tp:0 /drp:1
  //: joint g20 (w1) @(258, 636) /w:[ 2 -1 4 1 ]
  //: joint g15 (w4) @(265, 487) /w:[ 2 -1 4 1 ]
  //: joint g31 (clk) @(39, 524) /w:[ 10 12 -1 9 ]
  //: joint g29 (clk) @(39, 366) /w:[ 18 20 -1 17 ]
  //: IN g25 (clk) @(39,78) /sn:0 /R:3 /w:[ 33 ]
  //: OUT g17 (out) @(482,335) /sn:0 /w:[ 1 ]
  //: joint g14 (w6) @(258, 409) /w:[ 2 -1 4 1 ]
  FFD g5 (.D(w6), .Clk(clk), .Y(w4));   //: @(170, 468) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>11 Ro0<5 ]
  //: IN g21 (ctrlNeg) @(590,69) /sn:0 /R:2 /w:[ 0 ]
  //: joint g26 (clk) @(39, 109) /w:[ 30 32 -1 29 ]
  FFD g0 (.D(in), .Clk(clk), .Y(w2));   //: @(173, 50) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>31 Ro0<3 ]
  //: joint g22 (w2) @(262, 69) /w:[ 1 -1 2 4 ]
  FFD g18 (.D(w1), .Clk(clk), .Y(w0));   //: @(171, 708) /sz:(40, 40) /sn:0 /p:[ Li0>0 Bi0>0 Ro0<0 ]
  //: joint g12 (w9) @(256, 240) /w:[ 2 -1 4 1 ]
  //: joint g30 (clk) @(39, 448) /w:[ 14 16 -1 13 ]

endmodule
//: /netlistEnd

